`include "pulseChannel1.v"
`include "mixer.v"

`define PERIOD 4194304/16
`define LENGTH 10'd1023
`define PLAYBACK_LENGTH 10'd80
`define LONGREG reg [`LENGTH:0]

module gameboy();


	reg [31:0] [3:0] waveTable;

	// Square 1
	`LONGREG [2:0] sq1_swpPd;
	`LONGREG sq1_negate;
	`LONGREG [2:0] sq1_shift;
	`LONGREG [1:0] sq1_duty;
	`LONGREG [5:0] sq1_lenLoad;
	`LONGREG [3:0] sq1_startVol;
	`LONGREG sq1_envAdd;
	`LONGREG [2:0] sq1_period;
	`LONGREG [10:0] sq1_freq;
	`LONGREG sq1_trigger;
	`LONGREG sq1_lenEnable;

	`LONGREG [1:0] sq2_duty;
	`LONGREG [5:0] sq2_lenLoad;
	`LONGREG [3:0] sq2_startVol;
	`LONGREG sq2_envAdd;
	`LONGREG [2:0] sq2_period;
	`LONGREG [10:0] sq2_freq;
	`LONGREG sq2_trigger;
	`LONGREG sq2_lenEnable;

	wire clk; baseClk baseclk(clk);
	wire clk256; fixedTimer #(16384) tmr256(clk, clk256);
	wire clk128; fixedTimer #(2) tmr128(clk256, clk128);
	wire clk64; fixedTimer #(2) tmr64(clk128, clk64);

	wire clkT; fixedTimer #(`PERIOD) tmrT(clk, clkT);
	reg [$clog2(`LENGTH)-1:0] t;
	always @(posedge clkT) begin
		trigger = sq1_trigger[t];
		if (t < `PLAYBACK_LENGTH) t += 1;
		else $finish;
	end

	wire [3:0] sq1_out, sq2_out;
	reg trigger;

	pulseChannel1 pc1(clk, clk256, clk128, clk64, sq1_swpPd[t], sq1_negate[t], sq1_shift[t], sq1_freq[t], sq1_lenLoad[t], sq1_duty[t], sq1_startVol[t], sq1_period[t], sq1_lenEnable[t], trigger, sq1_envAdd[t], sq1_out);
	pulseChannel2 pc2(clk, clk256, clk128, clk64, sq2_freq[t], sq2_lenLoad[t], sq2_duty[t], sq2_startVol[t], sq2_period[t], sq2_lenEnable[t], trigger, sq2_envAdd[t], sq2_out);

	// Clock at falling edge so that nothing else is going on at the same time
	// swDac dac(!clk, sq1_out, sq2_out);
	mixer mxr(clk, 4'b1100, 4'b1100, 3'b111, 3'b111, sq1_out, sq2_out, 0, 0);

	reg [4:0] ii; // Fill in the wave table with a triangle wave

	initial begin
		t = 0;

		for (ii = 0; ii < 16; ii++) waveTable[ii] = {ii[3:0]};
		for (ii = 0; ii < 16; ii++) waveTable[ii+5'd16] = 4'd0 - {ii[3:0]};

sq1_swpPd[0] = 0.0;
 sq1_swpPd[1] = 0.0;
 sq1_swpPd[2] = 0.0;
 sq1_swpPd[3] = 0.0;
 sq1_swpPd[4] = 0.0;
 sq1_swpPd[5] = 0.0;
 sq1_swpPd[6] = 0.0;
 sq1_swpPd[7] = 0.0;
 sq1_swpPd[8] = 0.0;
 sq1_swpPd[9] = 0.0;
 sq1_swpPd[10] = 0.0;
 sq1_swpPd[11] = 0.0;
 sq1_swpPd[12] = 0.0;
 sq1_swpPd[13] = 0.0;
 sq1_swpPd[14] = 0.0;
 sq1_swpPd[15] = 0.0;
 sq1_swpPd[16] = 0.0;
 sq1_swpPd[17] = 0.0;
 sq1_swpPd[18] = 0.0;
 sq1_swpPd[19] = 0.0;
 sq1_swpPd[20] = 0.0;
 sq1_swpPd[21] = 0.0;
 sq1_swpPd[22] = 0.0;
 sq1_swpPd[23] = 0.0;
 sq1_swpPd[24] = 0.0;
 sq1_swpPd[25] = 0.0;
 sq1_swpPd[26] = 0.0;
 sq1_swpPd[27] = 0.0;
 sq1_swpPd[28] = 0.0;
 sq1_swpPd[29] = 0.0;
 sq1_swpPd[30] = 0.0;
 sq1_swpPd[31] = 0.0;
 sq1_swpPd[32] = 0.0;
 sq1_swpPd[33] = 0.0;
 sq1_swpPd[34] = 0.0;
 sq1_swpPd[35] = 0.0;
 sq1_swpPd[36] = 0.0;
 sq1_swpPd[37] = 0.0;
 sq1_swpPd[38] = 0.0;
 sq1_swpPd[39] = 0.0;
 sq1_swpPd[40] = 0.0;
 sq1_swpPd[41] = 0.0;
 sq1_swpPd[42] = 0.0;
 sq1_swpPd[43] = 0.0;
 sq1_swpPd[44] = 0.0;
 sq1_swpPd[45] = 0.0;
 sq1_swpPd[46] = 0.0;
 sq1_swpPd[47] = 0.0;
 sq1_swpPd[48] = 0.0;
 sq1_swpPd[49] = 0.0;
 sq1_swpPd[50] = 0.0;
 sq1_swpPd[51] = 0.0;
 sq1_swpPd[52] = 0.0;
 sq1_swpPd[53] = 0.0;
 sq1_swpPd[54] = 0.0;
 sq1_swpPd[55] = 0.0;
 sq1_swpPd[56] = 0.0;
 sq1_swpPd[57] = 0.0;
 sq1_swpPd[58] = 0.0;
 sq1_swpPd[59] = 0.0;
 sq1_swpPd[60] = 0.0;
 sq1_swpPd[61] = 0.0;
 sq1_swpPd[62] = 0.0;
 sq1_swpPd[63] = 0.0;
 sq1_swpPd[64] = 0.0;
 sq1_swpPd[65] = 0.0;
 sq1_swpPd[66] = 0.0;
 sq1_swpPd[67] = 0.0;
 sq1_swpPd[68] = 0.0;
 sq1_swpPd[69] = 0.0;
 sq1_swpPd[70] = 0.0;
 sq1_swpPd[71] = 0.0;
 sq1_swpPd[72] = 0.0;
 sq1_swpPd[73] = 0.0;
 sq1_swpPd[74] = 0.0;
 sq1_swpPd[75] = 0.0;
 sq1_swpPd[76] = 0.0;
 sq1_swpPd[77] = 0.0;
 sq1_swpPd[78] = 0.0;
 sq1_swpPd[79] = 0.0;
 sq1_swpPd[80] = 0.0;
 sq1_swpPd[81] = 0.0;
 sq1_swpPd[82] = 0.0;
 sq1_swpPd[83] = 0.0;
 sq1_swpPd[84] = 0.0;
 sq1_swpPd[85] = 0.0;
 sq1_swpPd[86] = 0.0;
 sq1_swpPd[87] = 0.0;
 sq1_swpPd[88] = 0.0;
 sq1_swpPd[89] = 0.0;
 sq1_swpPd[90] = 0.0;
 sq1_swpPd[91] = 0.0;
 sq1_swpPd[92] = 0.0;
 sq1_swpPd[93] = 0.0;
 sq1_swpPd[94] = 0.0;
 sq1_swpPd[95] = 0.0;
 sq1_swpPd[96] = 0.0;
 sq1_swpPd[97] = 0.0;
 sq1_swpPd[98] = 0.0;
 sq1_swpPd[99] = 0.0;
 sq1_swpPd[100] = 0.0;
 sq1_swpPd[101] = 0.0;
 sq1_swpPd[102] = 0.0;
 sq1_swpPd[103] = 0.0;
 sq1_swpPd[104] = 0.0;
 sq1_swpPd[105] = 0.0;
 sq1_swpPd[106] = 0.0;
 sq1_swpPd[107] = 0.0;
 sq1_swpPd[108] = 0.0;
 sq1_swpPd[109] = 0.0;
 sq1_swpPd[110] = 0.0;
 sq1_swpPd[111] = 0.0;
 sq1_swpPd[112] = 0.0;
 sq1_swpPd[113] = 0.0;
 sq1_swpPd[114] = 0.0;
 sq1_swpPd[115] = 0.0;
 sq1_swpPd[116] = 0.0;
 sq1_swpPd[117] = 0.0;
 sq1_swpPd[118] = 0.0;
 sq1_swpPd[119] = 0.0;
 sq1_swpPd[120] = 0.0;
 sq1_swpPd[121] = 0.0;
 sq1_swpPd[122] = 0.0;
 sq1_swpPd[123] = 0.0;
 sq1_swpPd[124] = 0.0;
 sq1_swpPd[125] = 0.0;
 sq1_swpPd[126] = 0.0;
 sq1_swpPd[127] = 0.0;
 sq1_swpPd[128] = 0.0;
 sq1_swpPd[129] = 0.0;
 sq1_swpPd[130] = 0.0;
 sq1_swpPd[131] = 0.0;
 sq1_swpPd[132] = 0.0;
 sq1_swpPd[133] = 0.0;
 sq1_swpPd[134] = 0.0;
 sq1_swpPd[135] = 0.0;
 sq1_swpPd[136] = 0.0;
 sq1_swpPd[137] = 0.0;
 sq1_swpPd[138] = 0.0;
 sq1_swpPd[139] = 0.0;
 sq1_swpPd[140] = 0.0;
 sq1_swpPd[141] = 0.0;
 sq1_swpPd[142] = 0.0;
 sq1_swpPd[143] = 0.0;
 sq1_swpPd[144] = 0.0;
 sq1_swpPd[145] = 0.0;
 sq1_swpPd[146] = 0.0;
 sq1_swpPd[147] = 0.0;
 sq1_swpPd[148] = 0.0;
 sq1_swpPd[149] = 0.0;
 sq1_swpPd[150] = 0.0;
 sq1_swpPd[151] = 0.0;
 sq1_swpPd[152] = 0.0;
 sq1_swpPd[153] = 0.0;
 sq1_swpPd[154] = 0.0;
 sq1_swpPd[155] = 0.0;
 sq1_swpPd[156] = 0.0;
 sq1_swpPd[157] = 0.0;
 sq1_swpPd[158] = 0.0;
 sq1_swpPd[159] = 0.0;
 sq1_swpPd[160] = 0.0;
 sq1_swpPd[161] = 0.0;
 sq1_swpPd[162] = 0.0;
 sq1_swpPd[163] = 0.0;
 sq1_swpPd[164] = 0.0;
 sq1_swpPd[165] = 0.0;
 sq1_swpPd[166] = 0.0;
 sq1_swpPd[167] = 0.0;
 sq1_swpPd[168] = 0.0;
 sq1_swpPd[169] = 0.0;
 sq1_swpPd[170] = 0.0;
 sq1_swpPd[171] = 0.0;
 sq1_swpPd[172] = 0.0;
 sq1_swpPd[173] = 0.0;
 sq1_swpPd[174] = 0.0;
 sq1_swpPd[175] = 0.0;
 sq1_swpPd[176] = 0.0;
 sq1_swpPd[177] = 0.0;
 sq1_swpPd[178] = 0.0;
 sq1_swpPd[179] = 0.0;
 sq1_swpPd[180] = 0.0;
 sq1_swpPd[181] = 0.0;
 sq1_swpPd[182] = 0.0;
 sq1_swpPd[183] = 0.0;
 sq1_swpPd[184] = 0.0;
 sq1_swpPd[185] = 0.0;
 sq1_swpPd[186] = 0.0;
 sq1_swpPd[187] = 0.0;
 sq1_swpPd[188] = 0.0;
 sq1_swpPd[189] = 0.0;
 sq1_swpPd[190] = 0.0;
 sq1_swpPd[191] = 0.0;
 sq1_swpPd[192] = 0.0;
 sq1_swpPd[193] = 0.0;
 sq1_swpPd[194] = 0.0;
 sq1_swpPd[195] = 0.0;
 sq1_swpPd[196] = 0.0;
 sq1_swpPd[197] = 0.0;
 sq1_swpPd[198] = 0.0;
 sq1_swpPd[199] = 0.0;
 sq1_swpPd[200] = 0.0;
 sq1_swpPd[201] = 0.0;
 sq1_swpPd[202] = 0.0;
 sq1_swpPd[203] = 0.0;
 sq1_swpPd[204] = 0.0;
 sq1_swpPd[205] = 0.0;
 sq1_swpPd[206] = 0.0;
 sq1_swpPd[207] = 0.0;
 sq1_swpPd[208] = 0.0;
 sq1_swpPd[209] = 0.0;
 sq1_swpPd[210] = 0.0;
 sq1_swpPd[211] = 0.0;
 sq1_swpPd[212] = 0.0;
 sq1_swpPd[213] = 0.0;
 sq1_swpPd[214] = 0.0;
 sq1_swpPd[215] = 0.0;
 sq1_swpPd[216] = 0.0;
 sq1_swpPd[217] = 0.0;
 sq1_swpPd[218] = 0.0;
 sq1_swpPd[219] = 0.0;
 sq1_swpPd[220] = 0.0;
 sq1_swpPd[221] = 0.0;
 sq1_swpPd[222] = 0.0;
 sq1_swpPd[223] = 0.0;
 sq1_swpPd[224] = 0.0;
 sq1_swpPd[225] = 0.0;
 sq1_swpPd[226] = 0.0;
 sq1_swpPd[227] = 0.0;
 sq1_swpPd[228] = 0.0;
 sq1_swpPd[229] = 0.0;
 sq1_swpPd[230] = 0.0;
 sq1_swpPd[231] = 0.0;
 sq1_swpPd[232] = 0.0;
 sq1_swpPd[233] = 0.0;
 sq1_swpPd[234] = 0.0;
 sq1_swpPd[235] = 0.0;
 sq1_swpPd[236] = 0.0;
 sq1_swpPd[237] = 0.0;
 sq1_swpPd[238] = 0.0;
 sq1_swpPd[239] = 0.0;
 sq1_swpPd[240] = 0.0;
 sq1_swpPd[241] = 0.0;
 sq1_swpPd[242] = 0.0;
 sq1_swpPd[243] = 0.0;
 sq1_swpPd[244] = 0.0;
 sq1_swpPd[245] = 0.0;
 sq1_swpPd[246] = 0.0;
 sq1_swpPd[247] = 0.0;
 sq1_swpPd[248] = 0.0;
 sq1_swpPd[249] = 0.0;
 sq1_swpPd[250] = 0.0;
 sq1_swpPd[251] = 0.0;
 sq1_swpPd[252] = 0.0;
 sq1_swpPd[253] = 0.0;
 sq1_swpPd[254] = 0.0;
 sq1_swpPd[255] = 0.0;
 sq1_swpPd[256] = 0.0;
 sq1_swpPd[257] = 0.0;
 sq1_swpPd[258] = 0.0;
 sq1_swpPd[259] = 0.0;
 sq1_swpPd[260] = 0.0;
 sq1_swpPd[261] = 0.0;
 sq1_swpPd[262] = 0.0;
 sq1_swpPd[263] = 0.0;
 sq1_swpPd[264] = 0.0;
 sq1_swpPd[265] = 0.0;
 sq1_swpPd[266] = 0.0;
 sq1_swpPd[267] = 0.0;
 sq1_swpPd[268] = 0.0;
 sq1_swpPd[269] = 0.0;
 sq1_swpPd[270] = 0.0;
 sq1_swpPd[271] = 0.0;
 sq1_swpPd[272] = 0.0;
 sq1_swpPd[273] = 0.0;
 sq1_swpPd[274] = 0.0;
 sq1_swpPd[275] = 0.0;
 sq1_swpPd[276] = 0.0;
 sq1_swpPd[277] = 0.0;
 sq1_swpPd[278] = 0.0;
 sq1_swpPd[279] = 0.0;
 sq1_swpPd[280] = 0.0;
 sq1_swpPd[281] = 0.0;
 sq1_swpPd[282] = 0.0;
 sq1_swpPd[283] = 0.0;
 sq1_swpPd[284] = 0.0;
 sq1_swpPd[285] = 0.0;
 sq1_swpPd[286] = 0.0;
 sq1_swpPd[287] = 0.0;
 sq1_swpPd[288] = 0.0;
 sq1_swpPd[289] = 0.0;
 sq1_swpPd[290] = 0.0;
 sq1_swpPd[291] = 0.0;
 sq1_swpPd[292] = 0.0;
 sq1_swpPd[293] = 0.0;
 sq1_swpPd[294] = 0.0;
 sq1_swpPd[295] = 0.0;
 sq1_swpPd[296] = 0.0;
 sq1_swpPd[297] = 0.0;
 sq1_swpPd[298] = 0.0;
 sq1_swpPd[299] = 0.0;
 sq1_swpPd[300] = 0.0;
 sq1_swpPd[301] = 0.0;
 sq1_swpPd[302] = 0.0;
 sq1_swpPd[303] = 0.0;
 sq1_swpPd[304] = 0.0;
 sq1_swpPd[305] = 0.0;
 sq1_swpPd[306] = 0.0;
 sq1_swpPd[307] = 0.0;
 sq1_swpPd[308] = 0.0;
 sq1_swpPd[309] = 0.0;
 sq1_swpPd[310] = 0.0;
 sq1_swpPd[311] = 0.0;
 sq1_swpPd[312] = 0.0;
 sq1_swpPd[313] = 0.0;
 sq1_swpPd[314] = 0.0;
 sq1_swpPd[315] = 0.0;
 sq1_swpPd[316] = 0.0;
 sq1_swpPd[317] = 0.0;
 sq1_swpPd[318] = 0.0;
 sq1_swpPd[319] = 0.0;
 sq1_swpPd[320] = 0.0;
 sq1_swpPd[321] = 0.0;
 sq1_swpPd[322] = 0.0;
 sq1_swpPd[323] = 0.0;
 sq1_swpPd[324] = 0.0;
 sq1_swpPd[325] = 0.0;
 sq1_swpPd[326] = 0.0;
 sq1_swpPd[327] = 0.0;
 sq1_swpPd[328] = 0.0;
 sq1_swpPd[329] = 0.0;
 sq1_swpPd[330] = 0.0;
 sq1_swpPd[331] = 0.0;
 sq1_swpPd[332] = 0.0;
 sq1_swpPd[333] = 0.0;
 sq1_swpPd[334] = 0.0;
 sq1_swpPd[335] = 0.0;
 sq1_swpPd[336] = 0.0;
 sq1_swpPd[337] = 0.0;
 sq1_swpPd[338] = 0.0;
 sq1_swpPd[339] = 0.0;
 sq1_swpPd[340] = 0.0;
 sq1_swpPd[341] = 0.0;
 sq1_swpPd[342] = 0.0;
 sq1_swpPd[343] = 0.0;
 sq1_swpPd[344] = 0.0;
 sq1_swpPd[345] = 0.0;
 sq1_swpPd[346] = 0.0;
 sq1_swpPd[347] = 0.0;
 sq1_swpPd[348] = 0.0;
 sq1_swpPd[349] = 0.0;
 sq1_swpPd[350] = 0.0;
 sq1_swpPd[351] = 0.0;
 sq1_swpPd[352] = 0.0;
 sq1_swpPd[353] = 0.0;
 sq1_swpPd[354] = 0.0;
 sq1_swpPd[355] = 0.0;
 sq1_swpPd[356] = 0.0;
 sq1_swpPd[357] = 0.0;
 sq1_swpPd[358] = 0.0;
 sq1_swpPd[359] = 0.0;
 sq1_swpPd[360] = 0.0;
 sq1_swpPd[361] = 0.0;
 sq1_swpPd[362] = 0.0;
 sq1_swpPd[363] = 0.0;
 sq1_swpPd[364] = 0.0;
 sq1_swpPd[365] = 0.0;
 sq1_swpPd[366] = 0.0;
 sq1_swpPd[367] = 0.0;
 sq1_swpPd[368] = 0.0;
 sq1_swpPd[369] = 0.0;
 sq1_swpPd[370] = 0.0;
 sq1_swpPd[371] = 0.0;
 sq1_swpPd[372] = 0.0;
 sq1_swpPd[373] = 0.0;
 sq1_swpPd[374] = 0.0;
 sq1_swpPd[375] = 0.0;
 sq1_swpPd[376] = 0.0;
 sq1_swpPd[377] = 0.0;
 sq1_swpPd[378] = 0.0;
 sq1_negate[0] = 0.0;
 sq1_negate[1] = 0.0;
 sq1_negate[2] = 0.0;
 sq1_negate[3] = 0.0;
 sq1_negate[4] = 0.0;
 sq1_negate[5] = 0.0;
 sq1_negate[6] = 0.0;
 sq1_negate[7] = 0.0;
 sq1_negate[8] = 0.0;
 sq1_negate[9] = 0.0;
 sq1_negate[10] = 0.0;
 sq1_negate[11] = 0.0;
 sq1_negate[12] = 0.0;
 sq1_negate[13] = 0.0;
 sq1_negate[14] = 0.0;
 sq1_negate[15] = 0.0;
 sq1_negate[16] = 0.0;
 sq1_negate[17] = 0.0;
 sq1_negate[18] = 0.0;
 sq1_negate[19] = 0.0;
 sq1_negate[20] = 0.0;
 sq1_negate[21] = 0.0;
 sq1_negate[22] = 0.0;
 sq1_negate[23] = 0.0;
 sq1_negate[24] = 0.0;
 sq1_negate[25] = 0.0;
 sq1_negate[26] = 0.0;
 sq1_negate[27] = 0.0;
 sq1_negate[28] = 0.0;
 sq1_negate[29] = 0.0;
 sq1_negate[30] = 0.0;
 sq1_negate[31] = 0.0;
 sq1_negate[32] = 0.0;
 sq1_negate[33] = 0.0;
 sq1_negate[34] = 0.0;
 sq1_negate[35] = 0.0;
 sq1_negate[36] = 0.0;
 sq1_negate[37] = 0.0;
 sq1_negate[38] = 0.0;
 sq1_negate[39] = 0.0;
 sq1_negate[40] = 0.0;
 sq1_negate[41] = 0.0;
 sq1_negate[42] = 0.0;
 sq1_negate[43] = 0.0;
 sq1_negate[44] = 0.0;
 sq1_negate[45] = 0.0;
 sq1_negate[46] = 0.0;
 sq1_negate[47] = 0.0;
 sq1_negate[48] = 0.0;
 sq1_negate[49] = 0.0;
 sq1_negate[50] = 0.0;
 sq1_negate[51] = 0.0;
 sq1_negate[52] = 0.0;
 sq1_negate[53] = 0.0;
 sq1_negate[54] = 0.0;
 sq1_negate[55] = 0.0;
 sq1_negate[56] = 0.0;
 sq1_negate[57] = 0.0;
 sq1_negate[58] = 0.0;
 sq1_negate[59] = 0.0;
 sq1_negate[60] = 0.0;
 sq1_negate[61] = 0.0;
 sq1_negate[62] = 0.0;
 sq1_negate[63] = 0.0;
 sq1_negate[64] = 0.0;
 sq1_negate[65] = 0.0;
 sq1_negate[66] = 0.0;
 sq1_negate[67] = 0.0;
 sq1_negate[68] = 0.0;
 sq1_negate[69] = 0.0;
 sq1_negate[70] = 0.0;
 sq1_negate[71] = 0.0;
 sq1_negate[72] = 0.0;
 sq1_negate[73] = 0.0;
 sq1_negate[74] = 0.0;
 sq1_negate[75] = 0.0;
 sq1_negate[76] = 0.0;
 sq1_negate[77] = 0.0;
 sq1_negate[78] = 0.0;
 sq1_negate[79] = 0.0;
 sq1_negate[80] = 0.0;
 sq1_negate[81] = 0.0;
 sq1_negate[82] = 0.0;
 sq1_negate[83] = 0.0;
 sq1_negate[84] = 0.0;
 sq1_negate[85] = 0.0;
 sq1_negate[86] = 0.0;
 sq1_negate[87] = 0.0;
 sq1_negate[88] = 0.0;
 sq1_negate[89] = 0.0;
 sq1_negate[90] = 0.0;
 sq1_negate[91] = 0.0;
 sq1_negate[92] = 0.0;
 sq1_negate[93] = 0.0;
 sq1_negate[94] = 0.0;
 sq1_negate[95] = 0.0;
 sq1_negate[96] = 0.0;
 sq1_negate[97] = 0.0;
 sq1_negate[98] = 0.0;
 sq1_negate[99] = 0.0;
 sq1_negate[100] = 0.0;
 sq1_negate[101] = 0.0;
 sq1_negate[102] = 0.0;
 sq1_negate[103] = 0.0;
 sq1_negate[104] = 0.0;
 sq1_negate[105] = 0.0;
 sq1_negate[106] = 0.0;
 sq1_negate[107] = 0.0;
 sq1_negate[108] = 0.0;
 sq1_negate[109] = 0.0;
 sq1_negate[110] = 0.0;
 sq1_negate[111] = 0.0;
 sq1_negate[112] = 0.0;
 sq1_negate[113] = 0.0;
 sq1_negate[114] = 0.0;
 sq1_negate[115] = 0.0;
 sq1_negate[116] = 0.0;
 sq1_negate[117] = 0.0;
 sq1_negate[118] = 0.0;
 sq1_negate[119] = 0.0;
 sq1_negate[120] = 0.0;
 sq1_negate[121] = 0.0;
 sq1_negate[122] = 0.0;
 sq1_negate[123] = 0.0;
 sq1_negate[124] = 0.0;
 sq1_negate[125] = 0.0;
 sq1_negate[126] = 0.0;
 sq1_negate[127] = 0.0;
 sq1_negate[128] = 0.0;
 sq1_negate[129] = 0.0;
 sq1_negate[130] = 0.0;
 sq1_negate[131] = 0.0;
 sq1_negate[132] = 0.0;
 sq1_negate[133] = 0.0;
 sq1_negate[134] = 0.0;
 sq1_negate[135] = 0.0;
 sq1_negate[136] = 0.0;
 sq1_negate[137] = 0.0;
 sq1_negate[138] = 0.0;
 sq1_negate[139] = 0.0;
 sq1_negate[140] = 0.0;
 sq1_negate[141] = 0.0;
 sq1_negate[142] = 0.0;
 sq1_negate[143] = 0.0;
 sq1_negate[144] = 0.0;
 sq1_negate[145] = 0.0;
 sq1_negate[146] = 0.0;
 sq1_negate[147] = 0.0;
 sq1_negate[148] = 0.0;
 sq1_negate[149] = 0.0;
 sq1_negate[150] = 0.0;
 sq1_negate[151] = 0.0;
 sq1_negate[152] = 0.0;
 sq1_negate[153] = 0.0;
 sq1_negate[154] = 0.0;
 sq1_negate[155] = 0.0;
 sq1_negate[156] = 0.0;
 sq1_negate[157] = 0.0;
 sq1_negate[158] = 0.0;
 sq1_negate[159] = 0.0;
 sq1_negate[160] = 0.0;
 sq1_negate[161] = 0.0;
 sq1_negate[162] = 0.0;
 sq1_negate[163] = 0.0;
 sq1_negate[164] = 0.0;
 sq1_negate[165] = 0.0;
 sq1_negate[166] = 0.0;
 sq1_negate[167] = 0.0;
 sq1_negate[168] = 0.0;
 sq1_negate[169] = 0.0;
 sq1_negate[170] = 0.0;
 sq1_negate[171] = 0.0;
 sq1_negate[172] = 0.0;
 sq1_negate[173] = 0.0;
 sq1_negate[174] = 0.0;
 sq1_negate[175] = 0.0;
 sq1_negate[176] = 0.0;
 sq1_negate[177] = 0.0;
 sq1_negate[178] = 0.0;
 sq1_negate[179] = 0.0;
 sq1_negate[180] = 0.0;
 sq1_negate[181] = 0.0;
 sq1_negate[182] = 0.0;
 sq1_negate[183] = 0.0;
 sq1_negate[184] = 0.0;
 sq1_negate[185] = 0.0;
 sq1_negate[186] = 0.0;
 sq1_negate[187] = 0.0;
 sq1_negate[188] = 0.0;
 sq1_negate[189] = 0.0;
 sq1_negate[190] = 0.0;
 sq1_negate[191] = 0.0;
 sq1_negate[192] = 0.0;
 sq1_negate[193] = 0.0;
 sq1_negate[194] = 0.0;
 sq1_negate[195] = 0.0;
 sq1_negate[196] = 0.0;
 sq1_negate[197] = 0.0;
 sq1_negate[198] = 0.0;
 sq1_negate[199] = 0.0;
 sq1_negate[200] = 0.0;
 sq1_negate[201] = 0.0;
 sq1_negate[202] = 0.0;
 sq1_negate[203] = 0.0;
 sq1_negate[204] = 0.0;
 sq1_negate[205] = 0.0;
 sq1_negate[206] = 0.0;
 sq1_negate[207] = 0.0;
 sq1_negate[208] = 0.0;
 sq1_negate[209] = 0.0;
 sq1_negate[210] = 0.0;
 sq1_negate[211] = 0.0;
 sq1_negate[212] = 0.0;
 sq1_negate[213] = 0.0;
 sq1_negate[214] = 0.0;
 sq1_negate[215] = 0.0;
 sq1_negate[216] = 0.0;
 sq1_negate[217] = 0.0;
 sq1_negate[218] = 0.0;
 sq1_negate[219] = 0.0;
 sq1_negate[220] = 0.0;
 sq1_negate[221] = 0.0;
 sq1_negate[222] = 0.0;
 sq1_negate[223] = 0.0;
 sq1_negate[224] = 0.0;
 sq1_negate[225] = 0.0;
 sq1_negate[226] = 0.0;
 sq1_negate[227] = 0.0;
 sq1_negate[228] = 0.0;
 sq1_negate[229] = 0.0;
 sq1_negate[230] = 0.0;
 sq1_negate[231] = 0.0;
 sq1_negate[232] = 0.0;
 sq1_negate[233] = 0.0;
 sq1_negate[234] = 0.0;
 sq1_negate[235] = 0.0;
 sq1_negate[236] = 0.0;
 sq1_negate[237] = 0.0;
 sq1_negate[238] = 0.0;
 sq1_negate[239] = 0.0;
 sq1_negate[240] = 0.0;
 sq1_negate[241] = 0.0;
 sq1_negate[242] = 0.0;
 sq1_negate[243] = 0.0;
 sq1_negate[244] = 0.0;
 sq1_negate[245] = 0.0;
 sq1_negate[246] = 0.0;
 sq1_negate[247] = 0.0;
 sq1_negate[248] = 0.0;
 sq1_negate[249] = 0.0;
 sq1_negate[250] = 0.0;
 sq1_negate[251] = 0.0;
 sq1_negate[252] = 0.0;
 sq1_negate[253] = 0.0;
 sq1_negate[254] = 0.0;
 sq1_negate[255] = 0.0;
 sq1_negate[256] = 0.0;
 sq1_negate[257] = 0.0;
 sq1_negate[258] = 0.0;
 sq1_negate[259] = 0.0;
 sq1_negate[260] = 0.0;
 sq1_negate[261] = 0.0;
 sq1_negate[262] = 0.0;
 sq1_negate[263] = 0.0;
 sq1_negate[264] = 0.0;
 sq1_negate[265] = 0.0;
 sq1_negate[266] = 0.0;
 sq1_negate[267] = 0.0;
 sq1_negate[268] = 0.0;
 sq1_negate[269] = 0.0;
 sq1_negate[270] = 0.0;
 sq1_negate[271] = 0.0;
 sq1_negate[272] = 0.0;
 sq1_negate[273] = 0.0;
 sq1_negate[274] = 0.0;
 sq1_negate[275] = 0.0;
 sq1_negate[276] = 0.0;
 sq1_negate[277] = 0.0;
 sq1_negate[278] = 0.0;
 sq1_negate[279] = 0.0;
 sq1_negate[280] = 0.0;
 sq1_negate[281] = 0.0;
 sq1_negate[282] = 0.0;
 sq1_negate[283] = 0.0;
 sq1_negate[284] = 0.0;
 sq1_negate[285] = 0.0;
 sq1_negate[286] = 0.0;
 sq1_negate[287] = 0.0;
 sq1_negate[288] = 0.0;
 sq1_negate[289] = 0.0;
 sq1_negate[290] = 0.0;
 sq1_negate[291] = 0.0;
 sq1_negate[292] = 0.0;
 sq1_negate[293] = 0.0;
 sq1_negate[294] = 0.0;
 sq1_negate[295] = 0.0;
 sq1_negate[296] = 0.0;
 sq1_negate[297] = 0.0;
 sq1_negate[298] = 0.0;
 sq1_negate[299] = 0.0;
 sq1_negate[300] = 0.0;
 sq1_negate[301] = 0.0;
 sq1_negate[302] = 0.0;
 sq1_negate[303] = 0.0;
 sq1_negate[304] = 0.0;
 sq1_negate[305] = 0.0;
 sq1_negate[306] = 0.0;
 sq1_negate[307] = 0.0;
 sq1_negate[308] = 0.0;
 sq1_negate[309] = 0.0;
 sq1_negate[310] = 0.0;
 sq1_negate[311] = 0.0;
 sq1_negate[312] = 0.0;
 sq1_negate[313] = 0.0;
 sq1_negate[314] = 0.0;
 sq1_negate[315] = 0.0;
 sq1_negate[316] = 0.0;
 sq1_negate[317] = 0.0;
 sq1_negate[318] = 0.0;
 sq1_negate[319] = 0.0;
 sq1_negate[320] = 0.0;
 sq1_negate[321] = 0.0;
 sq1_negate[322] = 0.0;
 sq1_negate[323] = 0.0;
 sq1_negate[324] = 0.0;
 sq1_negate[325] = 0.0;
 sq1_negate[326] = 0.0;
 sq1_negate[327] = 0.0;
 sq1_negate[328] = 0.0;
 sq1_negate[329] = 0.0;
 sq1_negate[330] = 0.0;
 sq1_negate[331] = 0.0;
 sq1_negate[332] = 0.0;
 sq1_negate[333] = 0.0;
 sq1_negate[334] = 0.0;
 sq1_negate[335] = 0.0;
 sq1_negate[336] = 0.0;
 sq1_negate[337] = 0.0;
 sq1_negate[338] = 0.0;
 sq1_negate[339] = 0.0;
 sq1_negate[340] = 0.0;
 sq1_negate[341] = 0.0;
 sq1_negate[342] = 0.0;
 sq1_negate[343] = 0.0;
 sq1_negate[344] = 0.0;
 sq1_negate[345] = 0.0;
 sq1_negate[346] = 0.0;
 sq1_negate[347] = 0.0;
 sq1_negate[348] = 0.0;
 sq1_negate[349] = 0.0;
 sq1_negate[350] = 0.0;
 sq1_negate[351] = 0.0;
 sq1_negate[352] = 0.0;
 sq1_negate[353] = 0.0;
 sq1_negate[354] = 0.0;
 sq1_negate[355] = 0.0;
 sq1_negate[356] = 0.0;
 sq1_negate[357] = 0.0;
 sq1_negate[358] = 0.0;
 sq1_negate[359] = 0.0;
 sq1_negate[360] = 0.0;
 sq1_negate[361] = 0.0;
 sq1_negate[362] = 0.0;
 sq1_negate[363] = 0.0;
 sq1_negate[364] = 0.0;
 sq1_negate[365] = 0.0;
 sq1_negate[366] = 0.0;
 sq1_negate[367] = 0.0;
 sq1_negate[368] = 0.0;
 sq1_negate[369] = 0.0;
 sq1_negate[370] = 0.0;
 sq1_negate[371] = 0.0;
 sq1_negate[372] = 0.0;
 sq1_negate[373] = 0.0;
 sq1_negate[374] = 0.0;
 sq1_negate[375] = 0.0;
 sq1_negate[376] = 0.0;
 sq1_negate[377] = 0.0;
 sq1_negate[378] = 0.0;
 sq1_shift[0] = 0.0;
 sq1_shift[1] = 0.0;
 sq1_shift[2] = 0.0;
 sq1_shift[3] = 0.0;
 sq1_shift[4] = 0.0;
 sq1_shift[5] = 0.0;
 sq1_shift[6] = 0.0;
 sq1_shift[7] = 0.0;
 sq1_shift[8] = 0.0;
 sq1_shift[9] = 0.0;
 sq1_shift[10] = 0.0;
 sq1_shift[11] = 0.0;
 sq1_shift[12] = 0.0;
 sq1_shift[13] = 0.0;
 sq1_shift[14] = 0.0;
 sq1_shift[15] = 0.0;
 sq1_shift[16] = 0.0;
 sq1_shift[17] = 0.0;
 sq1_shift[18] = 0.0;
 sq1_shift[19] = 0.0;
 sq1_shift[20] = 0.0;
 sq1_shift[21] = 0.0;
 sq1_shift[22] = 0.0;
 sq1_shift[23] = 0.0;
 sq1_shift[24] = 0.0;
 sq1_shift[25] = 0.0;
 sq1_shift[26] = 0.0;
 sq1_shift[27] = 0.0;
 sq1_shift[28] = 0.0;
 sq1_shift[29] = 0.0;
 sq1_shift[30] = 0.0;
 sq1_shift[31] = 0.0;
 sq1_shift[32] = 0.0;
 sq1_shift[33] = 0.0;
 sq1_shift[34] = 0.0;
 sq1_shift[35] = 0.0;
 sq1_shift[36] = 0.0;
 sq1_shift[37] = 0.0;
 sq1_shift[38] = 0.0;
 sq1_shift[39] = 0.0;
 sq1_shift[40] = 0.0;
 sq1_shift[41] = 0.0;
 sq1_shift[42] = 0.0;
 sq1_shift[43] = 0.0;
 sq1_shift[44] = 0.0;
 sq1_shift[45] = 0.0;
 sq1_shift[46] = 0.0;
 sq1_shift[47] = 0.0;
 sq1_shift[48] = 0.0;
 sq1_shift[49] = 0.0;
 sq1_shift[50] = 0.0;
 sq1_shift[51] = 0.0;
 sq1_shift[52] = 0.0;
 sq1_shift[53] = 0.0;
 sq1_shift[54] = 0.0;
 sq1_shift[55] = 0.0;
 sq1_shift[56] = 0.0;
 sq1_shift[57] = 0.0;
 sq1_shift[58] = 0.0;
 sq1_shift[59] = 0.0;
 sq1_shift[60] = 0.0;
 sq1_shift[61] = 0.0;
 sq1_shift[62] = 0.0;
 sq1_shift[63] = 0.0;
 sq1_shift[64] = 0.0;
 sq1_shift[65] = 0.0;
 sq1_shift[66] = 0.0;
 sq1_shift[67] = 0.0;
 sq1_shift[68] = 0.0;
 sq1_shift[69] = 0.0;
 sq1_shift[70] = 0.0;
 sq1_shift[71] = 0.0;
 sq1_shift[72] = 0.0;
 sq1_shift[73] = 0.0;
 sq1_shift[74] = 0.0;
 sq1_shift[75] = 0.0;
 sq1_shift[76] = 0.0;
 sq1_shift[77] = 0.0;
 sq1_shift[78] = 0.0;
 sq1_shift[79] = 0.0;
 sq1_shift[80] = 0.0;
 sq1_shift[81] = 0.0;
 sq1_shift[82] = 0.0;
 sq1_shift[83] = 0.0;
 sq1_shift[84] = 0.0;
 sq1_shift[85] = 0.0;
 sq1_shift[86] = 0.0;
 sq1_shift[87] = 0.0;
 sq1_shift[88] = 0.0;
 sq1_shift[89] = 0.0;
 sq1_shift[90] = 0.0;
 sq1_shift[91] = 0.0;
 sq1_shift[92] = 0.0;
 sq1_shift[93] = 0.0;
 sq1_shift[94] = 0.0;
 sq1_shift[95] = 0.0;
 sq1_shift[96] = 0.0;
 sq1_shift[97] = 0.0;
 sq1_shift[98] = 0.0;
 sq1_shift[99] = 0.0;
 sq1_shift[100] = 0.0;
 sq1_shift[101] = 0.0;
 sq1_shift[102] = 0.0;
 sq1_shift[103] = 0.0;
 sq1_shift[104] = 0.0;
 sq1_shift[105] = 0.0;
 sq1_shift[106] = 0.0;
 sq1_shift[107] = 0.0;
 sq1_shift[108] = 0.0;
 sq1_shift[109] = 0.0;
 sq1_shift[110] = 0.0;
 sq1_shift[111] = 0.0;
 sq1_shift[112] = 0.0;
 sq1_shift[113] = 0.0;
 sq1_shift[114] = 0.0;
 sq1_shift[115] = 0.0;
 sq1_shift[116] = 0.0;
 sq1_shift[117] = 0.0;
 sq1_shift[118] = 0.0;
 sq1_shift[119] = 0.0;
 sq1_shift[120] = 0.0;
 sq1_shift[121] = 0.0;
 sq1_shift[122] = 0.0;
 sq1_shift[123] = 0.0;
 sq1_shift[124] = 0.0;
 sq1_shift[125] = 0.0;
 sq1_shift[126] = 0.0;
 sq1_shift[127] = 0.0;
 sq1_shift[128] = 0.0;
 sq1_shift[129] = 0.0;
 sq1_shift[130] = 0.0;
 sq1_shift[131] = 0.0;
 sq1_shift[132] = 0.0;
 sq1_shift[133] = 0.0;
 sq1_shift[134] = 0.0;
 sq1_shift[135] = 0.0;
 sq1_shift[136] = 0.0;
 sq1_shift[137] = 0.0;
 sq1_shift[138] = 0.0;
 sq1_shift[139] = 0.0;
 sq1_shift[140] = 0.0;
 sq1_shift[141] = 0.0;
 sq1_shift[142] = 0.0;
 sq1_shift[143] = 0.0;
 sq1_shift[144] = 0.0;
 sq1_shift[145] = 0.0;
 sq1_shift[146] = 0.0;
 sq1_shift[147] = 0.0;
 sq1_shift[148] = 0.0;
 sq1_shift[149] = 0.0;
 sq1_shift[150] = 0.0;
 sq1_shift[151] = 0.0;
 sq1_shift[152] = 0.0;
 sq1_shift[153] = 0.0;
 sq1_shift[154] = 0.0;
 sq1_shift[155] = 0.0;
 sq1_shift[156] = 0.0;
 sq1_shift[157] = 0.0;
 sq1_shift[158] = 0.0;
 sq1_shift[159] = 0.0;
 sq1_shift[160] = 0.0;
 sq1_shift[161] = 0.0;
 sq1_shift[162] = 0.0;
 sq1_shift[163] = 0.0;
 sq1_shift[164] = 0.0;
 sq1_shift[165] = 0.0;
 sq1_shift[166] = 0.0;
 sq1_shift[167] = 0.0;
 sq1_shift[168] = 0.0;
 sq1_shift[169] = 0.0;
 sq1_shift[170] = 0.0;
 sq1_shift[171] = 0.0;
 sq1_shift[172] = 0.0;
 sq1_shift[173] = 0.0;
 sq1_shift[174] = 0.0;
 sq1_shift[175] = 0.0;
 sq1_shift[176] = 0.0;
 sq1_shift[177] = 0.0;
 sq1_shift[178] = 0.0;
 sq1_shift[179] = 0.0;
 sq1_shift[180] = 0.0;
 sq1_shift[181] = 0.0;
 sq1_shift[182] = 0.0;
 sq1_shift[183] = 0.0;
 sq1_shift[184] = 0.0;
 sq1_shift[185] = 0.0;
 sq1_shift[186] = 0.0;
 sq1_shift[187] = 0.0;
 sq1_shift[188] = 0.0;
 sq1_shift[189] = 0.0;
 sq1_shift[190] = 0.0;
 sq1_shift[191] = 0.0;
 sq1_shift[192] = 0.0;
 sq1_shift[193] = 0.0;
 sq1_shift[194] = 0.0;
 sq1_shift[195] = 0.0;
 sq1_shift[196] = 0.0;
 sq1_shift[197] = 0.0;
 sq1_shift[198] = 0.0;
 sq1_shift[199] = 0.0;
 sq1_shift[200] = 0.0;
 sq1_shift[201] = 0.0;
 sq1_shift[202] = 0.0;
 sq1_shift[203] = 0.0;
 sq1_shift[204] = 0.0;
 sq1_shift[205] = 0.0;
 sq1_shift[206] = 0.0;
 sq1_shift[207] = 0.0;
 sq1_shift[208] = 0.0;
 sq1_shift[209] = 0.0;
 sq1_shift[210] = 0.0;
 sq1_shift[211] = 0.0;
 sq1_shift[212] = 0.0;
 sq1_shift[213] = 0.0;
 sq1_shift[214] = 0.0;
 sq1_shift[215] = 0.0;
 sq1_shift[216] = 0.0;
 sq1_shift[217] = 0.0;
 sq1_shift[218] = 0.0;
 sq1_shift[219] = 0.0;
 sq1_shift[220] = 0.0;
 sq1_shift[221] = 0.0;
 sq1_shift[222] = 0.0;
 sq1_shift[223] = 0.0;
 sq1_shift[224] = 0.0;
 sq1_shift[225] = 0.0;
 sq1_shift[226] = 0.0;
 sq1_shift[227] = 0.0;
 sq1_shift[228] = 0.0;
 sq1_shift[229] = 0.0;
 sq1_shift[230] = 0.0;
 sq1_shift[231] = 0.0;
 sq1_shift[232] = 0.0;
 sq1_shift[233] = 0.0;
 sq1_shift[234] = 0.0;
 sq1_shift[235] = 0.0;
 sq1_shift[236] = 0.0;
 sq1_shift[237] = 0.0;
 sq1_shift[238] = 0.0;
 sq1_shift[239] = 0.0;
 sq1_shift[240] = 0.0;
 sq1_shift[241] = 0.0;
 sq1_shift[242] = 0.0;
 sq1_shift[243] = 0.0;
 sq1_shift[244] = 0.0;
 sq1_shift[245] = 0.0;
 sq1_shift[246] = 0.0;
 sq1_shift[247] = 0.0;
 sq1_shift[248] = 0.0;
 sq1_shift[249] = 0.0;
 sq1_shift[250] = 0.0;
 sq1_shift[251] = 0.0;
 sq1_shift[252] = 0.0;
 sq1_shift[253] = 0.0;
 sq1_shift[254] = 0.0;
 sq1_shift[255] = 0.0;
 sq1_shift[256] = 0.0;
 sq1_shift[257] = 0.0;
 sq1_shift[258] = 0.0;
 sq1_shift[259] = 0.0;
 sq1_shift[260] = 0.0;
 sq1_shift[261] = 0.0;
 sq1_shift[262] = 0.0;
 sq1_shift[263] = 0.0;
 sq1_shift[264] = 0.0;
 sq1_shift[265] = 0.0;
 sq1_shift[266] = 0.0;
 sq1_shift[267] = 0.0;
 sq1_shift[268] = 0.0;
 sq1_shift[269] = 0.0;
 sq1_shift[270] = 0.0;
 sq1_shift[271] = 0.0;
 sq1_shift[272] = 0.0;
 sq1_shift[273] = 0.0;
 sq1_shift[274] = 0.0;
 sq1_shift[275] = 0.0;
 sq1_shift[276] = 0.0;
 sq1_shift[277] = 0.0;
 sq1_shift[278] = 0.0;
 sq1_shift[279] = 0.0;
 sq1_shift[280] = 0.0;
 sq1_shift[281] = 0.0;
 sq1_shift[282] = 0.0;
 sq1_shift[283] = 0.0;
 sq1_shift[284] = 0.0;
 sq1_shift[285] = 0.0;
 sq1_shift[286] = 0.0;
 sq1_shift[287] = 0.0;
 sq1_shift[288] = 0.0;
 sq1_shift[289] = 0.0;
 sq1_shift[290] = 0.0;
 sq1_shift[291] = 0.0;
 sq1_shift[292] = 0.0;
 sq1_shift[293] = 0.0;
 sq1_shift[294] = 0.0;
 sq1_shift[295] = 0.0;
 sq1_shift[296] = 0.0;
 sq1_shift[297] = 0.0;
 sq1_shift[298] = 0.0;
 sq1_shift[299] = 0.0;
 sq1_shift[300] = 0.0;
 sq1_shift[301] = 0.0;
 sq1_shift[302] = 0.0;
 sq1_shift[303] = 0.0;
 sq1_shift[304] = 0.0;
 sq1_shift[305] = 0.0;
 sq1_shift[306] = 0.0;
 sq1_shift[307] = 0.0;
 sq1_shift[308] = 0.0;
 sq1_shift[309] = 0.0;
 sq1_shift[310] = 0.0;
 sq1_shift[311] = 0.0;
 sq1_shift[312] = 0.0;
 sq1_shift[313] = 0.0;
 sq1_shift[314] = 0.0;
 sq1_shift[315] = 0.0;
 sq1_shift[316] = 0.0;
 sq1_shift[317] = 0.0;
 sq1_shift[318] = 0.0;
 sq1_shift[319] = 0.0;
 sq1_shift[320] = 0.0;
 sq1_shift[321] = 0.0;
 sq1_shift[322] = 0.0;
 sq1_shift[323] = 0.0;
 sq1_shift[324] = 0.0;
 sq1_shift[325] = 0.0;
 sq1_shift[326] = 0.0;
 sq1_shift[327] = 0.0;
 sq1_shift[328] = 0.0;
 sq1_shift[329] = 0.0;
 sq1_shift[330] = 0.0;
 sq1_shift[331] = 0.0;
 sq1_shift[332] = 0.0;
 sq1_shift[333] = 0.0;
 sq1_shift[334] = 0.0;
 sq1_shift[335] = 0.0;
 sq1_shift[336] = 0.0;
 sq1_shift[337] = 0.0;
 sq1_shift[338] = 0.0;
 sq1_shift[339] = 0.0;
 sq1_shift[340] = 0.0;
 sq1_shift[341] = 0.0;
 sq1_shift[342] = 0.0;
 sq1_shift[343] = 0.0;
 sq1_shift[344] = 0.0;
 sq1_shift[345] = 0.0;
 sq1_shift[346] = 0.0;
 sq1_shift[347] = 0.0;
 sq1_shift[348] = 0.0;
 sq1_shift[349] = 0.0;
 sq1_shift[350] = 0.0;
 sq1_shift[351] = 0.0;
 sq1_shift[352] = 0.0;
 sq1_shift[353] = 0.0;
 sq1_shift[354] = 0.0;
 sq1_shift[355] = 0.0;
 sq1_shift[356] = 0.0;
 sq1_shift[357] = 0.0;
 sq1_shift[358] = 0.0;
 sq1_shift[359] = 0.0;
 sq1_shift[360] = 0.0;
 sq1_shift[361] = 0.0;
 sq1_shift[362] = 0.0;
 sq1_shift[363] = 0.0;
 sq1_shift[364] = 0.0;
 sq1_shift[365] = 0.0;
 sq1_shift[366] = 0.0;
 sq1_shift[367] = 0.0;
 sq1_shift[368] = 0.0;
 sq1_shift[369] = 0.0;
 sq1_shift[370] = 0.0;
 sq1_shift[371] = 0.0;
 sq1_shift[372] = 0.0;
 sq1_shift[373] = 0.0;
 sq1_shift[374] = 0.0;
 sq1_shift[375] = 0.0;
 sq1_shift[376] = 0.0;
 sq1_shift[377] = 0.0;
 sq1_shift[378] = 0.0;
 sq1_duty[0] = 2.0;
 sq1_duty[1] = 2.0;
 sq1_duty[2] = 2.0;
 sq1_duty[3] = 2.0;
 sq1_duty[4] = 2.0;
 sq1_duty[5] = 2.0;
 sq1_duty[6] = 2.0;
 sq1_duty[7] = 2.0;
 sq1_duty[8] = 2.0;
 sq1_duty[9] = 2.0;
 sq1_duty[10] = 2.0;
 sq1_duty[11] = 2.0;
 sq1_duty[12] = 2.0;
 sq1_duty[13] = 2.0;
 sq1_duty[14] = 2.0;
 sq1_duty[15] = 2.0;
 sq1_duty[16] = 2.0;
 sq1_duty[17] = 2.0;
 sq1_duty[18] = 2.0;
 sq1_duty[19] = 2.0;
 sq1_duty[20] = 2.0;
 sq1_duty[21] = 2.0;
 sq1_duty[22] = 2.0;
 sq1_duty[23] = 2.0;
 sq1_duty[24] = 2.0;
 sq1_duty[25] = 2.0;
 sq1_duty[26] = 2.0;
 sq1_duty[27] = 2.0;
 sq1_duty[28] = 2.0;
 sq1_duty[29] = 2.0;
 sq1_duty[30] = 2.0;
 sq1_duty[31] = 2.0;
 sq1_duty[32] = 2.0;
 sq1_duty[33] = 2.0;
 sq1_duty[34] = 2.0;
 sq1_duty[35] = 2.0;
 sq1_duty[36] = 2.0;
 sq1_duty[37] = 2.0;
 sq1_duty[38] = 2.0;
 sq1_duty[39] = 2.0;
 sq1_duty[40] = 2.0;
 sq1_duty[41] = 2.0;
 sq1_duty[42] = 2.0;
 sq1_duty[43] = 2.0;
 sq1_duty[44] = 2.0;
 sq1_duty[45] = 2.0;
 sq1_duty[46] = 2.0;
 sq1_duty[47] = 2.0;
 sq1_duty[48] = 2.0;
 sq1_duty[49] = 2.0;
 sq1_duty[50] = 2.0;
 sq1_duty[51] = 2.0;
 sq1_duty[52] = 2.0;
 sq1_duty[53] = 2.0;
 sq1_duty[54] = 2.0;
 sq1_duty[55] = 2.0;
 sq1_duty[56] = 2.0;
 sq1_duty[57] = 2.0;
 sq1_duty[58] = 2.0;
 sq1_duty[59] = 2.0;
 sq1_duty[60] = 2.0;
 sq1_duty[61] = 2.0;
 sq1_duty[62] = 2.0;
 sq1_duty[63] = 2.0;
 sq1_duty[64] = 2.0;
 sq1_duty[65] = 2.0;
 sq1_duty[66] = 2.0;
 sq1_duty[67] = 2.0;
 sq1_duty[68] = 2.0;
 sq1_duty[69] = 2.0;
 sq1_duty[70] = 2.0;
 sq1_duty[71] = 2.0;
 sq1_duty[72] = 2.0;
 sq1_duty[73] = 2.0;
 sq1_duty[74] = 2.0;
 sq1_duty[75] = 2.0;
 sq1_duty[76] = 2.0;
 sq1_duty[77] = 2.0;
 sq1_duty[78] = 2.0;
 sq1_duty[79] = 2.0;
 sq1_duty[80] = 2.0;
 sq1_duty[81] = 2.0;
 sq1_duty[82] = 2.0;
 sq1_duty[83] = 2.0;
 sq1_duty[84] = 2.0;
 sq1_duty[85] = 2.0;
 sq1_duty[86] = 2.0;
 sq1_duty[87] = 2.0;
 sq1_duty[88] = 2.0;
 sq1_duty[89] = 2.0;
 sq1_duty[90] = 2.0;
 sq1_duty[91] = 2.0;
 sq1_duty[92] = 2.0;
 sq1_duty[93] = 2.0;
 sq1_duty[94] = 2.0;
 sq1_duty[95] = 2.0;
 sq1_duty[96] = 2.0;
 sq1_duty[97] = 2.0;
 sq1_duty[98] = 2.0;
 sq1_duty[99] = 2.0;
 sq1_duty[100] = 2.0;
 sq1_duty[101] = 2.0;
 sq1_duty[102] = 2.0;
 sq1_duty[103] = 2.0;
 sq1_duty[104] = 2.0;
 sq1_duty[105] = 2.0;
 sq1_duty[106] = 2.0;
 sq1_duty[107] = 2.0;
 sq1_duty[108] = 2.0;
 sq1_duty[109] = 2.0;
 sq1_duty[110] = 2.0;
 sq1_duty[111] = 2.0;
 sq1_duty[112] = 2.0;
 sq1_duty[113] = 2.0;
 sq1_duty[114] = 2.0;
 sq1_duty[115] = 2.0;
 sq1_duty[116] = 2.0;
 sq1_duty[117] = 2.0;
 sq1_duty[118] = 2.0;
 sq1_duty[119] = 2.0;
 sq1_duty[120] = 2.0;
 sq1_duty[121] = 2.0;
 sq1_duty[122] = 2.0;
 sq1_duty[123] = 2.0;
 sq1_duty[124] = 2.0;
 sq1_duty[125] = 2.0;
 sq1_duty[126] = 2.0;
 sq1_duty[127] = 2.0;
 sq1_duty[128] = 2.0;
 sq1_duty[129] = 2.0;
 sq1_duty[130] = 2.0;
 sq1_duty[131] = 2.0;
 sq1_duty[132] = 2.0;
 sq1_duty[133] = 2.0;
 sq1_duty[134] = 2.0;
 sq1_duty[135] = 2.0;
 sq1_duty[136] = 2.0;
 sq1_duty[137] = 2.0;
 sq1_duty[138] = 2.0;
 sq1_duty[139] = 2.0;
 sq1_duty[140] = 2.0;
 sq1_duty[141] = 2.0;
 sq1_duty[142] = 2.0;
 sq1_duty[143] = 2.0;
 sq1_duty[144] = 2.0;
 sq1_duty[145] = 2.0;
 sq1_duty[146] = 2.0;
 sq1_duty[147] = 2.0;
 sq1_duty[148] = 2.0;
 sq1_duty[149] = 2.0;
 sq1_duty[150] = 2.0;
 sq1_duty[151] = 2.0;
 sq1_duty[152] = 2.0;
 sq1_duty[153] = 2.0;
 sq1_duty[154] = 2.0;
 sq1_duty[155] = 2.0;
 sq1_duty[156] = 2.0;
 sq1_duty[157] = 2.0;
 sq1_duty[158] = 2.0;
 sq1_duty[159] = 2.0;
 sq1_duty[160] = 2.0;
 sq1_duty[161] = 2.0;
 sq1_duty[162] = 2.0;
 sq1_duty[163] = 2.0;
 sq1_duty[164] = 2.0;
 sq1_duty[165] = 2.0;
 sq1_duty[166] = 2.0;
 sq1_duty[167] = 2.0;
 sq1_duty[168] = 2.0;
 sq1_duty[169] = 2.0;
 sq1_duty[170] = 2.0;
 sq1_duty[171] = 2.0;
 sq1_duty[172] = 2.0;
 sq1_duty[173] = 2.0;
 sq1_duty[174] = 2.0;
 sq1_duty[175] = 2.0;
 sq1_duty[176] = 2.0;
 sq1_duty[177] = 2.0;
 sq1_duty[178] = 2.0;
 sq1_duty[179] = 2.0;
 sq1_duty[180] = 2.0;
 sq1_duty[181] = 2.0;
 sq1_duty[182] = 2.0;
 sq1_duty[183] = 2.0;
 sq1_duty[184] = 2.0;
 sq1_duty[185] = 2.0;
 sq1_duty[186] = 2.0;
 sq1_duty[187] = 2.0;
 sq1_duty[188] = 2.0;
 sq1_duty[189] = 2.0;
 sq1_duty[190] = 2.0;
 sq1_duty[191] = 2.0;
 sq1_duty[192] = 2.0;
 sq1_duty[193] = 2.0;
 sq1_duty[194] = 2.0;
 sq1_duty[195] = 2.0;
 sq1_duty[196] = 2.0;
 sq1_duty[197] = 2.0;
 sq1_duty[198] = 2.0;
 sq1_duty[199] = 2.0;
 sq1_duty[200] = 2.0;
 sq1_duty[201] = 2.0;
 sq1_duty[202] = 2.0;
 sq1_duty[203] = 2.0;
 sq1_duty[204] = 2.0;
 sq1_duty[205] = 2.0;
 sq1_duty[206] = 2.0;
 sq1_duty[207] = 2.0;
 sq1_duty[208] = 2.0;
 sq1_duty[209] = 2.0;
 sq1_duty[210] = 2.0;
 sq1_duty[211] = 2.0;
 sq1_duty[212] = 2.0;
 sq1_duty[213] = 2.0;
 sq1_duty[214] = 2.0;
 sq1_duty[215] = 2.0;
 sq1_duty[216] = 2.0;
 sq1_duty[217] = 2.0;
 sq1_duty[218] = 2.0;
 sq1_duty[219] = 2.0;
 sq1_duty[220] = 2.0;
 sq1_duty[221] = 2.0;
 sq1_duty[222] = 2.0;
 sq1_duty[223] = 2.0;
 sq1_duty[224] = 2.0;
 sq1_duty[225] = 2.0;
 sq1_duty[226] = 2.0;
 sq1_duty[227] = 2.0;
 sq1_duty[228] = 2.0;
 sq1_duty[229] = 2.0;
 sq1_duty[230] = 2.0;
 sq1_duty[231] = 2.0;
 sq1_duty[232] = 2.0;
 sq1_duty[233] = 2.0;
 sq1_duty[234] = 2.0;
 sq1_duty[235] = 2.0;
 sq1_duty[236] = 2.0;
 sq1_duty[237] = 2.0;
 sq1_duty[238] = 2.0;
 sq1_duty[239] = 2.0;
 sq1_duty[240] = 2.0;
 sq1_duty[241] = 2.0;
 sq1_duty[242] = 2.0;
 sq1_duty[243] = 2.0;
 sq1_duty[244] = 2.0;
 sq1_duty[245] = 2.0;
 sq1_duty[246] = 2.0;
 sq1_duty[247] = 2.0;
 sq1_duty[248] = 2.0;
 sq1_duty[249] = 2.0;
 sq1_duty[250] = 2.0;
 sq1_duty[251] = 2.0;
 sq1_duty[252] = 2.0;
 sq1_duty[253] = 2.0;
 sq1_duty[254] = 2.0;
 sq1_duty[255] = 2.0;
 sq1_duty[256] = 2.0;
 sq1_duty[257] = 2.0;
 sq1_duty[258] = 2.0;
 sq1_duty[259] = 2.0;
 sq1_duty[260] = 2.0;
 sq1_duty[261] = 2.0;
 sq1_duty[262] = 2.0;
 sq1_duty[263] = 2.0;
 sq1_duty[264] = 2.0;
 sq1_duty[265] = 2.0;
 sq1_duty[266] = 2.0;
 sq1_duty[267] = 2.0;
 sq1_duty[268] = 2.0;
 sq1_duty[269] = 2.0;
 sq1_duty[270] = 2.0;
 sq1_duty[271] = 2.0;
 sq1_duty[272] = 2.0;
 sq1_duty[273] = 2.0;
 sq1_duty[274] = 2.0;
 sq1_duty[275] = 2.0;
 sq1_duty[276] = 2.0;
 sq1_duty[277] = 2.0;
 sq1_duty[278] = 2.0;
 sq1_duty[279] = 2.0;
 sq1_duty[280] = 2.0;
 sq1_duty[281] = 2.0;
 sq1_duty[282] = 2.0;
 sq1_duty[283] = 2.0;
 sq1_duty[284] = 2.0;
 sq1_duty[285] = 2.0;
 sq1_duty[286] = 2.0;
 sq1_duty[287] = 2.0;
 sq1_duty[288] = 2.0;
 sq1_duty[289] = 2.0;
 sq1_duty[290] = 2.0;
 sq1_duty[291] = 2.0;
 sq1_duty[292] = 2.0;
 sq1_duty[293] = 2.0;
 sq1_duty[294] = 2.0;
 sq1_duty[295] = 2.0;
 sq1_duty[296] = 2.0;
 sq1_duty[297] = 2.0;
 sq1_duty[298] = 2.0;
 sq1_duty[299] = 2.0;
 sq1_duty[300] = 2.0;
 sq1_duty[301] = 2.0;
 sq1_duty[302] = 2.0;
 sq1_duty[303] = 2.0;
 sq1_duty[304] = 2.0;
 sq1_duty[305] = 2.0;
 sq1_duty[306] = 2.0;
 sq1_duty[307] = 2.0;
 sq1_duty[308] = 2.0;
 sq1_duty[309] = 2.0;
 sq1_duty[310] = 2.0;
 sq1_duty[311] = 2.0;
 sq1_duty[312] = 2.0;
 sq1_duty[313] = 2.0;
 sq1_duty[314] = 2.0;
 sq1_duty[315] = 2.0;
 sq1_duty[316] = 2.0;
 sq1_duty[317] = 2.0;
 sq1_duty[318] = 2.0;
 sq1_duty[319] = 2.0;
 sq1_duty[320] = 2.0;
 sq1_duty[321] = 2.0;
 sq1_duty[322] = 2.0;
 sq1_duty[323] = 2.0;
 sq1_duty[324] = 2.0;
 sq1_duty[325] = 2.0;
 sq1_duty[326] = 2.0;
 sq1_duty[327] = 2.0;
 sq1_duty[328] = 2.0;
 sq1_duty[329] = 2.0;
 sq1_duty[330] = 2.0;
 sq1_duty[331] = 2.0;
 sq1_duty[332] = 2.0;
 sq1_duty[333] = 2.0;
 sq1_duty[334] = 2.0;
 sq1_duty[335] = 2.0;
 sq1_duty[336] = 2.0;
 sq1_duty[337] = 2.0;
 sq1_duty[338] = 2.0;
 sq1_duty[339] = 2.0;
 sq1_duty[340] = 2.0;
 sq1_duty[341] = 2.0;
 sq1_duty[342] = 2.0;
 sq1_duty[343] = 2.0;
 sq1_duty[344] = 2.0;
 sq1_duty[345] = 2.0;
 sq1_duty[346] = 2.0;
 sq1_duty[347] = 2.0;
 sq1_duty[348] = 2.0;
 sq1_duty[349] = 2.0;
 sq1_duty[350] = 2.0;
 sq1_duty[351] = 2.0;
 sq1_duty[352] = 2.0;
 sq1_duty[353] = 2.0;
 sq1_duty[354] = 2.0;
 sq1_duty[355] = 2.0;
 sq1_duty[356] = 2.0;
 sq1_duty[357] = 2.0;
 sq1_duty[358] = 2.0;
 sq1_duty[359] = 2.0;
 sq1_duty[360] = 2.0;
 sq1_duty[361] = 2.0;
 sq1_duty[362] = 2.0;
 sq1_duty[363] = 2.0;
 sq1_duty[364] = 2.0;
 sq1_duty[365] = 2.0;
 sq1_duty[366] = 2.0;
 sq1_duty[367] = 2.0;
 sq1_duty[368] = 2.0;
 sq1_duty[369] = 2.0;
 sq1_duty[370] = 2.0;
 sq1_duty[371] = 2.0;
 sq1_duty[372] = 2.0;
 sq1_duty[373] = 2.0;
 sq1_duty[374] = 2.0;
 sq1_duty[375] = 2.0;
 sq1_duty[376] = 2.0;
 sq1_duty[377] = 2.0;
 sq1_duty[378] = 2.0;
 sq1_lenLoad[0] = 32.0;
 sq1_lenLoad[1] = 32.0;
 sq1_lenLoad[2] = 32.0;
 sq1_lenLoad[3] = 32.0;
 sq1_lenLoad[4] = 32.0;
 sq1_lenLoad[5] = 32.0;
 sq1_lenLoad[6] = 32.0;
 sq1_lenLoad[7] = 32.0;
 sq1_lenLoad[8] = 32.0;
 sq1_lenLoad[9] = 32.0;
 sq1_lenLoad[10] = 32.0;
 sq1_lenLoad[11] = 32.0;
 sq1_lenLoad[12] = 32.0;
 sq1_lenLoad[13] = 32.0;
 sq1_lenLoad[14] = 32.0;
 sq1_lenLoad[15] = 32.0;
 sq1_lenLoad[16] = 32.0;
 sq1_lenLoad[17] = 32.0;
 sq1_lenLoad[18] = 32.0;
 sq1_lenLoad[19] = 32.0;
 sq1_lenLoad[20] = 32.0;
 sq1_lenLoad[21] = 32.0;
 sq1_lenLoad[22] = 32.0;
 sq1_lenLoad[23] = 32.0;
 sq1_lenLoad[24] = 32.0;
 sq1_lenLoad[25] = 32.0;
 sq1_lenLoad[26] = 32.0;
 sq1_lenLoad[27] = 32.0;
 sq1_lenLoad[28] = 32.0;
 sq1_lenLoad[29] = 32.0;
 sq1_lenLoad[30] = 32.0;
 sq1_lenLoad[31] = 32.0;
 sq1_lenLoad[32] = 32.0;
 sq1_lenLoad[33] = 32.0;
 sq1_lenLoad[34] = 32.0;
 sq1_lenLoad[35] = 32.0;
 sq1_lenLoad[36] = 32.0;
 sq1_lenLoad[37] = 32.0;
 sq1_lenLoad[38] = 32.0;
 sq1_lenLoad[39] = 32.0;
 sq1_lenLoad[40] = 32.0;
 sq1_lenLoad[41] = 32.0;
 sq1_lenLoad[42] = 32.0;
 sq1_lenLoad[43] = 32.0;
 sq1_lenLoad[44] = 32.0;
 sq1_lenLoad[45] = 32.0;
 sq1_lenLoad[46] = 32.0;
 sq1_lenLoad[47] = 32.0;
 sq1_lenLoad[48] = 32.0;
 sq1_lenLoad[49] = 32.0;
 sq1_lenLoad[50] = 32.0;
 sq1_lenLoad[51] = 32.0;
 sq1_lenLoad[52] = 32.0;
 sq1_lenLoad[53] = 32.0;
 sq1_lenLoad[54] = 32.0;
 sq1_lenLoad[55] = 32.0;
 sq1_lenLoad[56] = 32.0;
 sq1_lenLoad[57] = 32.0;
 sq1_lenLoad[58] = 32.0;
 sq1_lenLoad[59] = 32.0;
 sq1_lenLoad[60] = 32.0;
 sq1_lenLoad[61] = 32.0;
 sq1_lenLoad[62] = 32.0;
 sq1_lenLoad[63] = 32.0;
 sq1_lenLoad[64] = 32.0;
 sq1_lenLoad[65] = 32.0;
 sq1_lenLoad[66] = 32.0;
 sq1_lenLoad[67] = 32.0;
 sq1_lenLoad[68] = 32.0;
 sq1_lenLoad[69] = 32.0;
 sq1_lenLoad[70] = 32.0;
 sq1_lenLoad[71] = 32.0;
 sq1_lenLoad[72] = 32.0;
 sq1_lenLoad[73] = 32.0;
 sq1_lenLoad[74] = 32.0;
 sq1_lenLoad[75] = 32.0;
 sq1_lenLoad[76] = 32.0;
 sq1_lenLoad[77] = 32.0;
 sq1_lenLoad[78] = 32.0;
 sq1_lenLoad[79] = 32.0;
 sq1_lenLoad[80] = 32.0;
 sq1_lenLoad[81] = 32.0;
 sq1_lenLoad[82] = 32.0;
 sq1_lenLoad[83] = 32.0;
 sq1_lenLoad[84] = 32.0;
 sq1_lenLoad[85] = 32.0;
 sq1_lenLoad[86] = 32.0;
 sq1_lenLoad[87] = 32.0;
 sq1_lenLoad[88] = 32.0;
 sq1_lenLoad[89] = 32.0;
 sq1_lenLoad[90] = 32.0;
 sq1_lenLoad[91] = 32.0;
 sq1_lenLoad[92] = 32.0;
 sq1_lenLoad[93] = 32.0;
 sq1_lenLoad[94] = 32.0;
 sq1_lenLoad[95] = 32.0;
 sq1_lenLoad[96] = 32.0;
 sq1_lenLoad[97] = 32.0;
 sq1_lenLoad[98] = 32.0;
 sq1_lenLoad[99] = 32.0;
 sq1_lenLoad[100] = 32.0;
 sq1_lenLoad[101] = 32.0;
 sq1_lenLoad[102] = 32.0;
 sq1_lenLoad[103] = 32.0;
 sq1_lenLoad[104] = 32.0;
 sq1_lenLoad[105] = 32.0;
 sq1_lenLoad[106] = 32.0;
 sq1_lenLoad[107] = 32.0;
 sq1_lenLoad[108] = 32.0;
 sq1_lenLoad[109] = 32.0;
 sq1_lenLoad[110] = 32.0;
 sq1_lenLoad[111] = 32.0;
 sq1_lenLoad[112] = 32.0;
 sq1_lenLoad[113] = 32.0;
 sq1_lenLoad[114] = 32.0;
 sq1_lenLoad[115] = 32.0;
 sq1_lenLoad[116] = 32.0;
 sq1_lenLoad[117] = 32.0;
 sq1_lenLoad[118] = 32.0;
 sq1_lenLoad[119] = 32.0;
 sq1_lenLoad[120] = 32.0;
 sq1_lenLoad[121] = 32.0;
 sq1_lenLoad[122] = 32.0;
 sq1_lenLoad[123] = 32.0;
 sq1_lenLoad[124] = 32.0;
 sq1_lenLoad[125] = 32.0;
 sq1_lenLoad[126] = 32.0;
 sq1_lenLoad[127] = 32.0;
 sq1_lenLoad[128] = 32.0;
 sq1_lenLoad[129] = 32.0;
 sq1_lenLoad[130] = 32.0;
 sq1_lenLoad[131] = 32.0;
 sq1_lenLoad[132] = 32.0;
 sq1_lenLoad[133] = 32.0;
 sq1_lenLoad[134] = 32.0;
 sq1_lenLoad[135] = 32.0;
 sq1_lenLoad[136] = 32.0;
 sq1_lenLoad[137] = 32.0;
 sq1_lenLoad[138] = 32.0;
 sq1_lenLoad[139] = 32.0;
 sq1_lenLoad[140] = 32.0;
 sq1_lenLoad[141] = 32.0;
 sq1_lenLoad[142] = 32.0;
 sq1_lenLoad[143] = 32.0;
 sq1_lenLoad[144] = 32.0;
 sq1_lenLoad[145] = 32.0;
 sq1_lenLoad[146] = 32.0;
 sq1_lenLoad[147] = 32.0;
 sq1_lenLoad[148] = 32.0;
 sq1_lenLoad[149] = 32.0;
 sq1_lenLoad[150] = 32.0;
 sq1_lenLoad[151] = 32.0;
 sq1_lenLoad[152] = 32.0;
 sq1_lenLoad[153] = 32.0;
 sq1_lenLoad[154] = 32.0;
 sq1_lenLoad[155] = 32.0;
 sq1_lenLoad[156] = 32.0;
 sq1_lenLoad[157] = 32.0;
 sq1_lenLoad[158] = 32.0;
 sq1_lenLoad[159] = 32.0;
 sq1_lenLoad[160] = 32.0;
 sq1_lenLoad[161] = 32.0;
 sq1_lenLoad[162] = 32.0;
 sq1_lenLoad[163] = 32.0;
 sq1_lenLoad[164] = 32.0;
 sq1_lenLoad[165] = 32.0;
 sq1_lenLoad[166] = 32.0;
 sq1_lenLoad[167] = 32.0;
 sq1_lenLoad[168] = 32.0;
 sq1_lenLoad[169] = 32.0;
 sq1_lenLoad[170] = 32.0;
 sq1_lenLoad[171] = 32.0;
 sq1_lenLoad[172] = 32.0;
 sq1_lenLoad[173] = 32.0;
 sq1_lenLoad[174] = 32.0;
 sq1_lenLoad[175] = 32.0;
 sq1_lenLoad[176] = 32.0;
 sq1_lenLoad[177] = 32.0;
 sq1_lenLoad[178] = 32.0;
 sq1_lenLoad[179] = 32.0;
 sq1_lenLoad[180] = 32.0;
 sq1_lenLoad[181] = 32.0;
 sq1_lenLoad[182] = 32.0;
 sq1_lenLoad[183] = 32.0;
 sq1_lenLoad[184] = 32.0;
 sq1_lenLoad[185] = 32.0;
 sq1_lenLoad[186] = 32.0;
 sq1_lenLoad[187] = 32.0;
 sq1_lenLoad[188] = 32.0;
 sq1_lenLoad[189] = 32.0;
 sq1_lenLoad[190] = 32.0;
 sq1_lenLoad[191] = 32.0;
 sq1_lenLoad[192] = 32.0;
 sq1_lenLoad[193] = 32.0;
 sq1_lenLoad[194] = 32.0;
 sq1_lenLoad[195] = 32.0;
 sq1_lenLoad[196] = 32.0;
 sq1_lenLoad[197] = 32.0;
 sq1_lenLoad[198] = 32.0;
 sq1_lenLoad[199] = 32.0;
 sq1_lenLoad[200] = 32.0;
 sq1_lenLoad[201] = 32.0;
 sq1_lenLoad[202] = 32.0;
 sq1_lenLoad[203] = 32.0;
 sq1_lenLoad[204] = 32.0;
 sq1_lenLoad[205] = 32.0;
 sq1_lenLoad[206] = 32.0;
 sq1_lenLoad[207] = 32.0;
 sq1_lenLoad[208] = 32.0;
 sq1_lenLoad[209] = 32.0;
 sq1_lenLoad[210] = 32.0;
 sq1_lenLoad[211] = 32.0;
 sq1_lenLoad[212] = 32.0;
 sq1_lenLoad[213] = 32.0;
 sq1_lenLoad[214] = 32.0;
 sq1_lenLoad[215] = 32.0;
 sq1_lenLoad[216] = 32.0;
 sq1_lenLoad[217] = 32.0;
 sq1_lenLoad[218] = 32.0;
 sq1_lenLoad[219] = 32.0;
 sq1_lenLoad[220] = 32.0;
 sq1_lenLoad[221] = 32.0;
 sq1_lenLoad[222] = 32.0;
 sq1_lenLoad[223] = 32.0;
 sq1_lenLoad[224] = 32.0;
 sq1_lenLoad[225] = 32.0;
 sq1_lenLoad[226] = 32.0;
 sq1_lenLoad[227] = 32.0;
 sq1_lenLoad[228] = 32.0;
 sq1_lenLoad[229] = 32.0;
 sq1_lenLoad[230] = 32.0;
 sq1_lenLoad[231] = 32.0;
 sq1_lenLoad[232] = 32.0;
 sq1_lenLoad[233] = 32.0;
 sq1_lenLoad[234] = 32.0;
 sq1_lenLoad[235] = 32.0;
 sq1_lenLoad[236] = 32.0;
 sq1_lenLoad[237] = 32.0;
 sq1_lenLoad[238] = 32.0;
 sq1_lenLoad[239] = 32.0;
 sq1_lenLoad[240] = 32.0;
 sq1_lenLoad[241] = 32.0;
 sq1_lenLoad[242] = 32.0;
 sq1_lenLoad[243] = 32.0;
 sq1_lenLoad[244] = 32.0;
 sq1_lenLoad[245] = 32.0;
 sq1_lenLoad[246] = 32.0;
 sq1_lenLoad[247] = 32.0;
 sq1_lenLoad[248] = 32.0;
 sq1_lenLoad[249] = 32.0;
 sq1_lenLoad[250] = 32.0;
 sq1_lenLoad[251] = 32.0;
 sq1_lenLoad[252] = 32.0;
 sq1_lenLoad[253] = 32.0;
 sq1_lenLoad[254] = 32.0;
 sq1_lenLoad[255] = 32.0;
 sq1_lenLoad[256] = 32.0;
 sq1_lenLoad[257] = 32.0;
 sq1_lenLoad[258] = 32.0;
 sq1_lenLoad[259] = 32.0;
 sq1_lenLoad[260] = 32.0;
 sq1_lenLoad[261] = 32.0;
 sq1_lenLoad[262] = 32.0;
 sq1_lenLoad[263] = 32.0;
 sq1_lenLoad[264] = 32.0;
 sq1_lenLoad[265] = 32.0;
 sq1_lenLoad[266] = 32.0;
 sq1_lenLoad[267] = 32.0;
 sq1_lenLoad[268] = 32.0;
 sq1_lenLoad[269] = 32.0;
 sq1_lenLoad[270] = 32.0;
 sq1_lenLoad[271] = 32.0;
 sq1_lenLoad[272] = 32.0;
 sq1_lenLoad[273] = 32.0;
 sq1_lenLoad[274] = 32.0;
 sq1_lenLoad[275] = 32.0;
 sq1_lenLoad[276] = 32.0;
 sq1_lenLoad[277] = 32.0;
 sq1_lenLoad[278] = 32.0;
 sq1_lenLoad[279] = 32.0;
 sq1_lenLoad[280] = 32.0;
 sq1_lenLoad[281] = 32.0;
 sq1_lenLoad[282] = 32.0;
 sq1_lenLoad[283] = 32.0;
 sq1_lenLoad[284] = 32.0;
 sq1_lenLoad[285] = 32.0;
 sq1_lenLoad[286] = 32.0;
 sq1_lenLoad[287] = 32.0;
 sq1_lenLoad[288] = 32.0;
 sq1_lenLoad[289] = 32.0;
 sq1_lenLoad[290] = 32.0;
 sq1_lenLoad[291] = 32.0;
 sq1_lenLoad[292] = 32.0;
 sq1_lenLoad[293] = 32.0;
 sq1_lenLoad[294] = 32.0;
 sq1_lenLoad[295] = 32.0;
 sq1_lenLoad[296] = 32.0;
 sq1_lenLoad[297] = 32.0;
 sq1_lenLoad[298] = 32.0;
 sq1_lenLoad[299] = 32.0;
 sq1_lenLoad[300] = 32.0;
 sq1_lenLoad[301] = 32.0;
 sq1_lenLoad[302] = 32.0;
 sq1_lenLoad[303] = 32.0;
 sq1_lenLoad[304] = 32.0;
 sq1_lenLoad[305] = 32.0;
 sq1_lenLoad[306] = 32.0;
 sq1_lenLoad[307] = 32.0;
 sq1_lenLoad[308] = 32.0;
 sq1_lenLoad[309] = 32.0;
 sq1_lenLoad[310] = 32.0;
 sq1_lenLoad[311] = 32.0;
 sq1_lenLoad[312] = 32.0;
 sq1_lenLoad[313] = 32.0;
 sq1_lenLoad[314] = 32.0;
 sq1_lenLoad[315] = 32.0;
 sq1_lenLoad[316] = 32.0;
 sq1_lenLoad[317] = 32.0;
 sq1_lenLoad[318] = 32.0;
 sq1_lenLoad[319] = 32.0;
 sq1_lenLoad[320] = 32.0;
 sq1_lenLoad[321] = 32.0;
 sq1_lenLoad[322] = 32.0;
 sq1_lenLoad[323] = 32.0;
 sq1_lenLoad[324] = 32.0;
 sq1_lenLoad[325] = 32.0;
 sq1_lenLoad[326] = 32.0;
 sq1_lenLoad[327] = 32.0;
 sq1_lenLoad[328] = 32.0;
 sq1_lenLoad[329] = 32.0;
 sq1_lenLoad[330] = 32.0;
 sq1_lenLoad[331] = 32.0;
 sq1_lenLoad[332] = 32.0;
 sq1_lenLoad[333] = 32.0;
 sq1_lenLoad[334] = 32.0;
 sq1_lenLoad[335] = 32.0;
 sq1_lenLoad[336] = 32.0;
 sq1_lenLoad[337] = 32.0;
 sq1_lenLoad[338] = 32.0;
 sq1_lenLoad[339] = 32.0;
 sq1_lenLoad[340] = 32.0;
 sq1_lenLoad[341] = 32.0;
 sq1_lenLoad[342] = 32.0;
 sq1_lenLoad[343] = 32.0;
 sq1_lenLoad[344] = 32.0;
 sq1_lenLoad[345] = 32.0;
 sq1_lenLoad[346] = 32.0;
 sq1_lenLoad[347] = 32.0;
 sq1_lenLoad[348] = 32.0;
 sq1_lenLoad[349] = 32.0;
 sq1_lenLoad[350] = 32.0;
 sq1_lenLoad[351] = 32.0;
 sq1_lenLoad[352] = 32.0;
 sq1_lenLoad[353] = 32.0;
 sq1_lenLoad[354] = 32.0;
 sq1_lenLoad[355] = 32.0;
 sq1_lenLoad[356] = 32.0;
 sq1_lenLoad[357] = 32.0;
 sq1_lenLoad[358] = 32.0;
 sq1_lenLoad[359] = 32.0;
 sq1_lenLoad[360] = 32.0;
 sq1_lenLoad[361] = 32.0;
 sq1_lenLoad[362] = 32.0;
 sq1_lenLoad[363] = 32.0;
 sq1_lenLoad[364] = 32.0;
 sq1_lenLoad[365] = 32.0;
 sq1_lenLoad[366] = 32.0;
 sq1_lenLoad[367] = 32.0;
 sq1_lenLoad[368] = 32.0;
 sq1_lenLoad[369] = 32.0;
 sq1_lenLoad[370] = 32.0;
 sq1_lenLoad[371] = 32.0;
 sq1_lenLoad[372] = 32.0;
 sq1_lenLoad[373] = 32.0;
 sq1_lenLoad[374] = 32.0;
 sq1_lenLoad[375] = 32.0;
 sq1_lenLoad[376] = 32.0;
 sq1_lenLoad[377] = 32.0;
 sq1_lenLoad[378] = 32.0;
 sq1_startVol[0] = 12.0;
 sq1_startVol[1] = 12.0;
 sq1_startVol[2] = 12.0;
 sq1_startVol[3] = 12.0;
 sq1_startVol[4] = 12.0;
 sq1_startVol[5] = 12.0;
 sq1_startVol[6] = 12.0;
 sq1_startVol[7] = 12.0;
 sq1_startVol[8] = 12.0;
 sq1_startVol[9] = 12.0;
 sq1_startVol[10] = 12.0;
 sq1_startVol[11] = 12.0;
 sq1_startVol[12] = 12.0;
 sq1_startVol[13] = 12.0;
 sq1_startVol[14] = 12.0;
 sq1_startVol[15] = 12.0;
 sq1_startVol[16] = 12.0;
 sq1_startVol[17] = 12.0;
 sq1_startVol[18] = 12.0;
 sq1_startVol[19] = 12.0;
 sq1_startVol[20] = 12.0;
 sq1_startVol[21] = 12.0;
 sq1_startVol[22] = 12.0;
 sq1_startVol[23] = 12.0;
 sq1_startVol[24] = 12.0;
 sq1_startVol[25] = 12.0;
 sq1_startVol[26] = 12.0;
 sq1_startVol[27] = 12.0;
 sq1_startVol[28] = 12.0;
 sq1_startVol[29] = 12.0;
 sq1_startVol[30] = 12.0;
 sq1_startVol[31] = 12.0;
 sq1_startVol[32] = 12.0;
 sq1_startVol[33] = 12.0;
 sq1_startVol[34] = 12.0;
 sq1_startVol[35] = 12.0;
 sq1_startVol[36] = 12.0;
 sq1_startVol[37] = 12.0;
 sq1_startVol[38] = 12.0;
 sq1_startVol[39] = 12.0;
 sq1_startVol[40] = 12.0;
 sq1_startVol[41] = 12.0;
 sq1_startVol[42] = 12.0;
 sq1_startVol[43] = 12.0;
 sq1_startVol[44] = 12.0;
 sq1_startVol[45] = 12.0;
 sq1_startVol[46] = 12.0;
 sq1_startVol[47] = 12.0;
 sq1_startVol[48] = 12.0;
 sq1_startVol[49] = 12.0;
 sq1_startVol[50] = 12.0;
 sq1_startVol[51] = 12.0;
 sq1_startVol[52] = 12.0;
 sq1_startVol[53] = 12.0;
 sq1_startVol[54] = 12.0;
 sq1_startVol[55] = 12.0;
 sq1_startVol[56] = 12.0;
 sq1_startVol[57] = 12.0;
 sq1_startVol[58] = 12.0;
 sq1_startVol[59] = 12.0;
 sq1_startVol[60] = 12.0;
 sq1_startVol[61] = 12.0;
 sq1_startVol[62] = 12.0;
 sq1_startVol[63] = 12.0;
 sq1_startVol[64] = 12.0;
 sq1_startVol[65] = 12.0;
 sq1_startVol[66] = 12.0;
 sq1_startVol[67] = 12.0;
 sq1_startVol[68] = 12.0;
 sq1_startVol[69] = 12.0;
 sq1_startVol[70] = 12.0;
 sq1_startVol[71] = 12.0;
 sq1_startVol[72] = 12.0;
 sq1_startVol[73] = 12.0;
 sq1_startVol[74] = 12.0;
 sq1_startVol[75] = 12.0;
 sq1_startVol[76] = 12.0;
 sq1_startVol[77] = 12.0;
 sq1_startVol[78] = 12.0;
 sq1_startVol[79] = 12.0;
 sq1_startVol[80] = 12.0;
 sq1_startVol[81] = 12.0;
 sq1_startVol[82] = 12.0;
 sq1_startVol[83] = 12.0;
 sq1_startVol[84] = 12.0;
 sq1_startVol[85] = 12.0;
 sq1_startVol[86] = 12.0;
 sq1_startVol[87] = 12.0;
 sq1_startVol[88] = 12.0;
 sq1_startVol[89] = 12.0;
 sq1_startVol[90] = 12.0;
 sq1_startVol[91] = 12.0;
 sq1_startVol[92] = 12.0;
 sq1_startVol[93] = 12.0;
 sq1_startVol[94] = 12.0;
 sq1_startVol[95] = 12.0;
 sq1_startVol[96] = 12.0;
 sq1_startVol[97] = 12.0;
 sq1_startVol[98] = 12.0;
 sq1_startVol[99] = 12.0;
 sq1_startVol[100] = 12.0;
 sq1_startVol[101] = 12.0;
 sq1_startVol[102] = 12.0;
 sq1_startVol[103] = 12.0;
 sq1_startVol[104] = 12.0;
 sq1_startVol[105] = 12.0;
 sq1_startVol[106] = 12.0;
 sq1_startVol[107] = 12.0;
 sq1_startVol[108] = 12.0;
 sq1_startVol[109] = 12.0;
 sq1_startVol[110] = 12.0;
 sq1_startVol[111] = 12.0;
 sq1_startVol[112] = 12.0;
 sq1_startVol[113] = 12.0;
 sq1_startVol[114] = 12.0;
 sq1_startVol[115] = 12.0;
 sq1_startVol[116] = 12.0;
 sq1_startVol[117] = 12.0;
 sq1_startVol[118] = 12.0;
 sq1_startVol[119] = 12.0;
 sq1_startVol[120] = 12.0;
 sq1_startVol[121] = 12.0;
 sq1_startVol[122] = 12.0;
 sq1_startVol[123] = 12.0;
 sq1_startVol[124] = 12.0;
 sq1_startVol[125] = 12.0;
 sq1_startVol[126] = 12.0;
 sq1_startVol[127] = 12.0;
 sq1_startVol[128] = 12.0;
 sq1_startVol[129] = 12.0;
 sq1_startVol[130] = 12.0;
 sq1_startVol[131] = 12.0;
 sq1_startVol[132] = 12.0;
 sq1_startVol[133] = 12.0;
 sq1_startVol[134] = 12.0;
 sq1_startVol[135] = 12.0;
 sq1_startVol[136] = 12.0;
 sq1_startVol[137] = 12.0;
 sq1_startVol[138] = 12.0;
 sq1_startVol[139] = 12.0;
 sq1_startVol[140] = 12.0;
 sq1_startVol[141] = 12.0;
 sq1_startVol[142] = 12.0;
 sq1_startVol[143] = 12.0;
 sq1_startVol[144] = 12.0;
 sq1_startVol[145] = 12.0;
 sq1_startVol[146] = 12.0;
 sq1_startVol[147] = 12.0;
 sq1_startVol[148] = 12.0;
 sq1_startVol[149] = 12.0;
 sq1_startVol[150] = 12.0;
 sq1_startVol[151] = 12.0;
 sq1_startVol[152] = 12.0;
 sq1_startVol[153] = 12.0;
 sq1_startVol[154] = 12.0;
 sq1_startVol[155] = 12.0;
 sq1_startVol[156] = 12.0;
 sq1_startVol[157] = 12.0;
 sq1_startVol[158] = 12.0;
 sq1_startVol[159] = 12.0;
 sq1_startVol[160] = 12.0;
 sq1_startVol[161] = 12.0;
 sq1_startVol[162] = 12.0;
 sq1_startVol[163] = 12.0;
 sq1_startVol[164] = 12.0;
 sq1_startVol[165] = 12.0;
 sq1_startVol[166] = 12.0;
 sq1_startVol[167] = 12.0;
 sq1_startVol[168] = 12.0;
 sq1_startVol[169] = 12.0;
 sq1_startVol[170] = 12.0;
 sq1_startVol[171] = 12.0;
 sq1_startVol[172] = 12.0;
 sq1_startVol[173] = 12.0;
 sq1_startVol[174] = 12.0;
 sq1_startVol[175] = 12.0;
 sq1_startVol[176] = 12.0;
 sq1_startVol[177] = 12.0;
 sq1_startVol[178] = 12.0;
 sq1_startVol[179] = 12.0;
 sq1_startVol[180] = 12.0;
 sq1_startVol[181] = 12.0;
 sq1_startVol[182] = 12.0;
 sq1_startVol[183] = 12.0;
 sq1_startVol[184] = 12.0;
 sq1_startVol[185] = 12.0;
 sq1_startVol[186] = 12.0;
 sq1_startVol[187] = 12.0;
 sq1_startVol[188] = 12.0;
 sq1_startVol[189] = 12.0;
 sq1_startVol[190] = 12.0;
 sq1_startVol[191] = 12.0;
 sq1_startVol[192] = 12.0;
 sq1_startVol[193] = 12.0;
 sq1_startVol[194] = 12.0;
 sq1_startVol[195] = 12.0;
 sq1_startVol[196] = 12.0;
 sq1_startVol[197] = 12.0;
 sq1_startVol[198] = 12.0;
 sq1_startVol[199] = 12.0;
 sq1_startVol[200] = 12.0;
 sq1_startVol[201] = 12.0;
 sq1_startVol[202] = 12.0;
 sq1_startVol[203] = 12.0;
 sq1_startVol[204] = 12.0;
 sq1_startVol[205] = 12.0;
 sq1_startVol[206] = 12.0;
 sq1_startVol[207] = 12.0;
 sq1_startVol[208] = 12.0;
 sq1_startVol[209] = 12.0;
 sq1_startVol[210] = 12.0;
 sq1_startVol[211] = 12.0;
 sq1_startVol[212] = 12.0;
 sq1_startVol[213] = 12.0;
 sq1_startVol[214] = 12.0;
 sq1_startVol[215] = 12.0;
 sq1_startVol[216] = 12.0;
 sq1_startVol[217] = 12.0;
 sq1_startVol[218] = 12.0;
 sq1_startVol[219] = 12.0;
 sq1_startVol[220] = 12.0;
 sq1_startVol[221] = 12.0;
 sq1_startVol[222] = 12.0;
 sq1_startVol[223] = 12.0;
 sq1_startVol[224] = 12.0;
 sq1_startVol[225] = 12.0;
 sq1_startVol[226] = 12.0;
 sq1_startVol[227] = 12.0;
 sq1_startVol[228] = 12.0;
 sq1_startVol[229] = 12.0;
 sq1_startVol[230] = 12.0;
 sq1_startVol[231] = 12.0;
 sq1_startVol[232] = 12.0;
 sq1_startVol[233] = 12.0;
 sq1_startVol[234] = 12.0;
 sq1_startVol[235] = 12.0;
 sq1_startVol[236] = 12.0;
 sq1_startVol[237] = 12.0;
 sq1_startVol[238] = 12.0;
 sq1_startVol[239] = 12.0;
 sq1_startVol[240] = 12.0;
 sq1_startVol[241] = 12.0;
 sq1_startVol[242] = 12.0;
 sq1_startVol[243] = 12.0;
 sq1_startVol[244] = 12.0;
 sq1_startVol[245] = 12.0;
 sq1_startVol[246] = 12.0;
 sq1_startVol[247] = 12.0;
 sq1_startVol[248] = 12.0;
 sq1_startVol[249] = 12.0;
 sq1_startVol[250] = 12.0;
 sq1_startVol[251] = 12.0;
 sq1_startVol[252] = 12.0;
 sq1_startVol[253] = 12.0;
 sq1_startVol[254] = 12.0;
 sq1_startVol[255] = 12.0;
 sq1_startVol[256] = 12.0;
 sq1_startVol[257] = 12.0;
 sq1_startVol[258] = 12.0;
 sq1_startVol[259] = 12.0;
 sq1_startVol[260] = 12.0;
 sq1_startVol[261] = 12.0;
 sq1_startVol[262] = 12.0;
 sq1_startVol[263] = 12.0;
 sq1_startVol[264] = 12.0;
 sq1_startVol[265] = 12.0;
 sq1_startVol[266] = 12.0;
 sq1_startVol[267] = 12.0;
 sq1_startVol[268] = 12.0;
 sq1_startVol[269] = 12.0;
 sq1_startVol[270] = 12.0;
 sq1_startVol[271] = 12.0;
 sq1_startVol[272] = 12.0;
 sq1_startVol[273] = 12.0;
 sq1_startVol[274] = 12.0;
 sq1_startVol[275] = 12.0;
 sq1_startVol[276] = 12.0;
 sq1_startVol[277] = 12.0;
 sq1_startVol[278] = 12.0;
 sq1_startVol[279] = 12.0;
 sq1_startVol[280] = 12.0;
 sq1_startVol[281] = 12.0;
 sq1_startVol[282] = 12.0;
 sq1_startVol[283] = 12.0;
 sq1_startVol[284] = 12.0;
 sq1_startVol[285] = 12.0;
 sq1_startVol[286] = 12.0;
 sq1_startVol[287] = 12.0;
 sq1_startVol[288] = 12.0;
 sq1_startVol[289] = 12.0;
 sq1_startVol[290] = 12.0;
 sq1_startVol[291] = 12.0;
 sq1_startVol[292] = 12.0;
 sq1_startVol[293] = 12.0;
 sq1_startVol[294] = 12.0;
 sq1_startVol[295] = 12.0;
 sq1_startVol[296] = 12.0;
 sq1_startVol[297] = 12.0;
 sq1_startVol[298] = 12.0;
 sq1_startVol[299] = 12.0;
 sq1_startVol[300] = 12.0;
 sq1_startVol[301] = 12.0;
 sq1_startVol[302] = 12.0;
 sq1_startVol[303] = 12.0;
 sq1_startVol[304] = 12.0;
 sq1_startVol[305] = 12.0;
 sq1_startVol[306] = 12.0;
 sq1_startVol[307] = 12.0;
 sq1_startVol[308] = 12.0;
 sq1_startVol[309] = 12.0;
 sq1_startVol[310] = 12.0;
 sq1_startVol[311] = 12.0;
 sq1_startVol[312] = 12.0;
 sq1_startVol[313] = 12.0;
 sq1_startVol[314] = 12.0;
 sq1_startVol[315] = 12.0;
 sq1_startVol[316] = 12.0;
 sq1_startVol[317] = 12.0;
 sq1_startVol[318] = 12.0;
 sq1_startVol[319] = 12.0;
 sq1_startVol[320] = 12.0;
 sq1_startVol[321] = 12.0;
 sq1_startVol[322] = 12.0;
 sq1_startVol[323] = 12.0;
 sq1_startVol[324] = 12.0;
 sq1_startVol[325] = 12.0;
 sq1_startVol[326] = 12.0;
 sq1_startVol[327] = 12.0;
 sq1_startVol[328] = 12.0;
 sq1_startVol[329] = 12.0;
 sq1_startVol[330] = 12.0;
 sq1_startVol[331] = 12.0;
 sq1_startVol[332] = 12.0;
 sq1_startVol[333] = 12.0;
 sq1_startVol[334] = 12.0;
 sq1_startVol[335] = 12.0;
 sq1_startVol[336] = 12.0;
 sq1_startVol[337] = 12.0;
 sq1_startVol[338] = 12.0;
 sq1_startVol[339] = 12.0;
 sq1_startVol[340] = 12.0;
 sq1_startVol[341] = 12.0;
 sq1_startVol[342] = 12.0;
 sq1_startVol[343] = 12.0;
 sq1_startVol[344] = 12.0;
 sq1_startVol[345] = 12.0;
 sq1_startVol[346] = 12.0;
 sq1_startVol[347] = 12.0;
 sq1_startVol[348] = 12.0;
 sq1_startVol[349] = 12.0;
 sq1_startVol[350] = 12.0;
 sq1_startVol[351] = 12.0;
 sq1_startVol[352] = 12.0;
 sq1_startVol[353] = 12.0;
 sq1_startVol[354] = 12.0;
 sq1_startVol[355] = 12.0;
 sq1_startVol[356] = 12.0;
 sq1_startVol[357] = 12.0;
 sq1_startVol[358] = 12.0;
 sq1_startVol[359] = 12.0;
 sq1_startVol[360] = 12.0;
 sq1_startVol[361] = 12.0;
 sq1_startVol[362] = 12.0;
 sq1_startVol[363] = 12.0;
 sq1_startVol[364] = 12.0;
 sq1_startVol[365] = 12.0;
 sq1_startVol[366] = 12.0;
 sq1_startVol[367] = 12.0;
 sq1_startVol[368] = 12.0;
 sq1_startVol[369] = 12.0;
 sq1_startVol[370] = 12.0;
 sq1_startVol[371] = 12.0;
 sq1_startVol[372] = 12.0;
 sq1_startVol[373] = 12.0;
 sq1_startVol[374] = 12.0;
 sq1_startVol[375] = 12.0;
 sq1_startVol[376] = 12.0;
 sq1_startVol[377] = 12.0;
 sq1_startVol[378] = 12.0;
 sq1_envAdd[0] = 0.0;
 sq1_envAdd[1] = 0.0;
 sq1_envAdd[2] = 0.0;
 sq1_envAdd[3] = 0.0;
 sq1_envAdd[4] = 0.0;
 sq1_envAdd[5] = 0.0;
 sq1_envAdd[6] = 0.0;
 sq1_envAdd[7] = 0.0;
 sq1_envAdd[8] = 0.0;
 sq1_envAdd[9] = 0.0;
 sq1_envAdd[10] = 0.0;
 sq1_envAdd[11] = 0.0;
 sq1_envAdd[12] = 0.0;
 sq1_envAdd[13] = 0.0;
 sq1_envAdd[14] = 0.0;
 sq1_envAdd[15] = 0.0;
 sq1_envAdd[16] = 0.0;
 sq1_envAdd[17] = 0.0;
 sq1_envAdd[18] = 0.0;
 sq1_envAdd[19] = 0.0;
 sq1_envAdd[20] = 0.0;
 sq1_envAdd[21] = 0.0;
 sq1_envAdd[22] = 0.0;
 sq1_envAdd[23] = 0.0;
 sq1_envAdd[24] = 0.0;
 sq1_envAdd[25] = 0.0;
 sq1_envAdd[26] = 0.0;
 sq1_envAdd[27] = 0.0;
 sq1_envAdd[28] = 0.0;
 sq1_envAdd[29] = 0.0;
 sq1_envAdd[30] = 0.0;
 sq1_envAdd[31] = 0.0;
 sq1_envAdd[32] = 0.0;
 sq1_envAdd[33] = 0.0;
 sq1_envAdd[34] = 0.0;
 sq1_envAdd[35] = 0.0;
 sq1_envAdd[36] = 0.0;
 sq1_envAdd[37] = 0.0;
 sq1_envAdd[38] = 0.0;
 sq1_envAdd[39] = 0.0;
 sq1_envAdd[40] = 0.0;
 sq1_envAdd[41] = 0.0;
 sq1_envAdd[42] = 0.0;
 sq1_envAdd[43] = 0.0;
 sq1_envAdd[44] = 0.0;
 sq1_envAdd[45] = 0.0;
 sq1_envAdd[46] = 0.0;
 sq1_envAdd[47] = 0.0;
 sq1_envAdd[48] = 0.0;
 sq1_envAdd[49] = 0.0;
 sq1_envAdd[50] = 0.0;
 sq1_envAdd[51] = 0.0;
 sq1_envAdd[52] = 0.0;
 sq1_envAdd[53] = 0.0;
 sq1_envAdd[54] = 0.0;
 sq1_envAdd[55] = 0.0;
 sq1_envAdd[56] = 0.0;
 sq1_envAdd[57] = 0.0;
 sq1_envAdd[58] = 0.0;
 sq1_envAdd[59] = 0.0;
 sq1_envAdd[60] = 0.0;
 sq1_envAdd[61] = 0.0;
 sq1_envAdd[62] = 0.0;
 sq1_envAdd[63] = 0.0;
 sq1_envAdd[64] = 0.0;
 sq1_envAdd[65] = 0.0;
 sq1_envAdd[66] = 0.0;
 sq1_envAdd[67] = 0.0;
 sq1_envAdd[68] = 0.0;
 sq1_envAdd[69] = 0.0;
 sq1_envAdd[70] = 0.0;
 sq1_envAdd[71] = 0.0;
 sq1_envAdd[72] = 0.0;
 sq1_envAdd[73] = 0.0;
 sq1_envAdd[74] = 0.0;
 sq1_envAdd[75] = 0.0;
 sq1_envAdd[76] = 0.0;
 sq1_envAdd[77] = 0.0;
 sq1_envAdd[78] = 0.0;
 sq1_envAdd[79] = 0.0;
 sq1_envAdd[80] = 0.0;
 sq1_envAdd[81] = 0.0;
 sq1_envAdd[82] = 0.0;
 sq1_envAdd[83] = 0.0;
 sq1_envAdd[84] = 0.0;
 sq1_envAdd[85] = 0.0;
 sq1_envAdd[86] = 0.0;
 sq1_envAdd[87] = 0.0;
 sq1_envAdd[88] = 0.0;
 sq1_envAdd[89] = 0.0;
 sq1_envAdd[90] = 0.0;
 sq1_envAdd[91] = 0.0;
 sq1_envAdd[92] = 0.0;
 sq1_envAdd[93] = 0.0;
 sq1_envAdd[94] = 0.0;
 sq1_envAdd[95] = 0.0;
 sq1_envAdd[96] = 0.0;
 sq1_envAdd[97] = 0.0;
 sq1_envAdd[98] = 0.0;
 sq1_envAdd[99] = 0.0;
 sq1_envAdd[100] = 0.0;
 sq1_envAdd[101] = 0.0;
 sq1_envAdd[102] = 0.0;
 sq1_envAdd[103] = 0.0;
 sq1_envAdd[104] = 0.0;
 sq1_envAdd[105] = 0.0;
 sq1_envAdd[106] = 0.0;
 sq1_envAdd[107] = 0.0;
 sq1_envAdd[108] = 0.0;
 sq1_envAdd[109] = 0.0;
 sq1_envAdd[110] = 0.0;
 sq1_envAdd[111] = 0.0;
 sq1_envAdd[112] = 0.0;
 sq1_envAdd[113] = 0.0;
 sq1_envAdd[114] = 0.0;
 sq1_envAdd[115] = 0.0;
 sq1_envAdd[116] = 0.0;
 sq1_envAdd[117] = 0.0;
 sq1_envAdd[118] = 0.0;
 sq1_envAdd[119] = 0.0;
 sq1_envAdd[120] = 0.0;
 sq1_envAdd[121] = 0.0;
 sq1_envAdd[122] = 0.0;
 sq1_envAdd[123] = 0.0;
 sq1_envAdd[124] = 0.0;
 sq1_envAdd[125] = 0.0;
 sq1_envAdd[126] = 0.0;
 sq1_envAdd[127] = 0.0;
 sq1_envAdd[128] = 0.0;
 sq1_envAdd[129] = 0.0;
 sq1_envAdd[130] = 0.0;
 sq1_envAdd[131] = 0.0;
 sq1_envAdd[132] = 0.0;
 sq1_envAdd[133] = 0.0;
 sq1_envAdd[134] = 0.0;
 sq1_envAdd[135] = 0.0;
 sq1_envAdd[136] = 0.0;
 sq1_envAdd[137] = 0.0;
 sq1_envAdd[138] = 0.0;
 sq1_envAdd[139] = 0.0;
 sq1_envAdd[140] = 0.0;
 sq1_envAdd[141] = 0.0;
 sq1_envAdd[142] = 0.0;
 sq1_envAdd[143] = 0.0;
 sq1_envAdd[144] = 0.0;
 sq1_envAdd[145] = 0.0;
 sq1_envAdd[146] = 0.0;
 sq1_envAdd[147] = 0.0;
 sq1_envAdd[148] = 0.0;
 sq1_envAdd[149] = 0.0;
 sq1_envAdd[150] = 0.0;
 sq1_envAdd[151] = 0.0;
 sq1_envAdd[152] = 0.0;
 sq1_envAdd[153] = 0.0;
 sq1_envAdd[154] = 0.0;
 sq1_envAdd[155] = 0.0;
 sq1_envAdd[156] = 0.0;
 sq1_envAdd[157] = 0.0;
 sq1_envAdd[158] = 0.0;
 sq1_envAdd[159] = 0.0;
 sq1_envAdd[160] = 0.0;
 sq1_envAdd[161] = 0.0;
 sq1_envAdd[162] = 0.0;
 sq1_envAdd[163] = 0.0;
 sq1_envAdd[164] = 0.0;
 sq1_envAdd[165] = 0.0;
 sq1_envAdd[166] = 0.0;
 sq1_envAdd[167] = 0.0;
 sq1_envAdd[168] = 0.0;
 sq1_envAdd[169] = 0.0;
 sq1_envAdd[170] = 0.0;
 sq1_envAdd[171] = 0.0;
 sq1_envAdd[172] = 0.0;
 sq1_envAdd[173] = 0.0;
 sq1_envAdd[174] = 0.0;
 sq1_envAdd[175] = 0.0;
 sq1_envAdd[176] = 0.0;
 sq1_envAdd[177] = 0.0;
 sq1_envAdd[178] = 0.0;
 sq1_envAdd[179] = 0.0;
 sq1_envAdd[180] = 0.0;
 sq1_envAdd[181] = 0.0;
 sq1_envAdd[182] = 0.0;
 sq1_envAdd[183] = 0.0;
 sq1_envAdd[184] = 0.0;
 sq1_envAdd[185] = 0.0;
 sq1_envAdd[186] = 0.0;
 sq1_envAdd[187] = 0.0;
 sq1_envAdd[188] = 0.0;
 sq1_envAdd[189] = 0.0;
 sq1_envAdd[190] = 0.0;
 sq1_envAdd[191] = 0.0;
 sq1_envAdd[192] = 0.0;
 sq1_envAdd[193] = 0.0;
 sq1_envAdd[194] = 0.0;
 sq1_envAdd[195] = 0.0;
 sq1_envAdd[196] = 0.0;
 sq1_envAdd[197] = 0.0;
 sq1_envAdd[198] = 0.0;
 sq1_envAdd[199] = 0.0;
 sq1_envAdd[200] = 0.0;
 sq1_envAdd[201] = 0.0;
 sq1_envAdd[202] = 0.0;
 sq1_envAdd[203] = 0.0;
 sq1_envAdd[204] = 0.0;
 sq1_envAdd[205] = 0.0;
 sq1_envAdd[206] = 0.0;
 sq1_envAdd[207] = 0.0;
 sq1_envAdd[208] = 0.0;
 sq1_envAdd[209] = 0.0;
 sq1_envAdd[210] = 0.0;
 sq1_envAdd[211] = 0.0;
 sq1_envAdd[212] = 0.0;
 sq1_envAdd[213] = 0.0;
 sq1_envAdd[214] = 0.0;
 sq1_envAdd[215] = 0.0;
 sq1_envAdd[216] = 0.0;
 sq1_envAdd[217] = 0.0;
 sq1_envAdd[218] = 0.0;
 sq1_envAdd[219] = 0.0;
 sq1_envAdd[220] = 0.0;
 sq1_envAdd[221] = 0.0;
 sq1_envAdd[222] = 0.0;
 sq1_envAdd[223] = 0.0;
 sq1_envAdd[224] = 0.0;
 sq1_envAdd[225] = 0.0;
 sq1_envAdd[226] = 0.0;
 sq1_envAdd[227] = 0.0;
 sq1_envAdd[228] = 0.0;
 sq1_envAdd[229] = 0.0;
 sq1_envAdd[230] = 0.0;
 sq1_envAdd[231] = 0.0;
 sq1_envAdd[232] = 0.0;
 sq1_envAdd[233] = 0.0;
 sq1_envAdd[234] = 0.0;
 sq1_envAdd[235] = 0.0;
 sq1_envAdd[236] = 0.0;
 sq1_envAdd[237] = 0.0;
 sq1_envAdd[238] = 0.0;
 sq1_envAdd[239] = 0.0;
 sq1_envAdd[240] = 0.0;
 sq1_envAdd[241] = 0.0;
 sq1_envAdd[242] = 0.0;
 sq1_envAdd[243] = 0.0;
 sq1_envAdd[244] = 0.0;
 sq1_envAdd[245] = 0.0;
 sq1_envAdd[246] = 0.0;
 sq1_envAdd[247] = 0.0;
 sq1_envAdd[248] = 0.0;
 sq1_envAdd[249] = 0.0;
 sq1_envAdd[250] = 0.0;
 sq1_envAdd[251] = 0.0;
 sq1_envAdd[252] = 0.0;
 sq1_envAdd[253] = 0.0;
 sq1_envAdd[254] = 0.0;
 sq1_envAdd[255] = 0.0;
 sq1_envAdd[256] = 0.0;
 sq1_envAdd[257] = 0.0;
 sq1_envAdd[258] = 0.0;
 sq1_envAdd[259] = 0.0;
 sq1_envAdd[260] = 0.0;
 sq1_envAdd[261] = 0.0;
 sq1_envAdd[262] = 0.0;
 sq1_envAdd[263] = 0.0;
 sq1_envAdd[264] = 0.0;
 sq1_envAdd[265] = 0.0;
 sq1_envAdd[266] = 0.0;
 sq1_envAdd[267] = 0.0;
 sq1_envAdd[268] = 0.0;
 sq1_envAdd[269] = 0.0;
 sq1_envAdd[270] = 0.0;
 sq1_envAdd[271] = 0.0;
 sq1_envAdd[272] = 0.0;
 sq1_envAdd[273] = 0.0;
 sq1_envAdd[274] = 0.0;
 sq1_envAdd[275] = 0.0;
 sq1_envAdd[276] = 0.0;
 sq1_envAdd[277] = 0.0;
 sq1_envAdd[278] = 0.0;
 sq1_envAdd[279] = 0.0;
 sq1_envAdd[280] = 0.0;
 sq1_envAdd[281] = 0.0;
 sq1_envAdd[282] = 0.0;
 sq1_envAdd[283] = 0.0;
 sq1_envAdd[284] = 0.0;
 sq1_envAdd[285] = 0.0;
 sq1_envAdd[286] = 0.0;
 sq1_envAdd[287] = 0.0;
 sq1_envAdd[288] = 0.0;
 sq1_envAdd[289] = 0.0;
 sq1_envAdd[290] = 0.0;
 sq1_envAdd[291] = 0.0;
 sq1_envAdd[292] = 0.0;
 sq1_envAdd[293] = 0.0;
 sq1_envAdd[294] = 0.0;
 sq1_envAdd[295] = 0.0;
 sq1_envAdd[296] = 0.0;
 sq1_envAdd[297] = 0.0;
 sq1_envAdd[298] = 0.0;
 sq1_envAdd[299] = 0.0;
 sq1_envAdd[300] = 0.0;
 sq1_envAdd[301] = 0.0;
 sq1_envAdd[302] = 0.0;
 sq1_envAdd[303] = 0.0;
 sq1_envAdd[304] = 0.0;
 sq1_envAdd[305] = 0.0;
 sq1_envAdd[306] = 0.0;
 sq1_envAdd[307] = 0.0;
 sq1_envAdd[308] = 0.0;
 sq1_envAdd[309] = 0.0;
 sq1_envAdd[310] = 0.0;
 sq1_envAdd[311] = 0.0;
 sq1_envAdd[312] = 0.0;
 sq1_envAdd[313] = 0.0;
 sq1_envAdd[314] = 0.0;
 sq1_envAdd[315] = 0.0;
 sq1_envAdd[316] = 0.0;
 sq1_envAdd[317] = 0.0;
 sq1_envAdd[318] = 0.0;
 sq1_envAdd[319] = 0.0;
 sq1_envAdd[320] = 0.0;
 sq1_envAdd[321] = 0.0;
 sq1_envAdd[322] = 0.0;
 sq1_envAdd[323] = 0.0;
 sq1_envAdd[324] = 0.0;
 sq1_envAdd[325] = 0.0;
 sq1_envAdd[326] = 0.0;
 sq1_envAdd[327] = 0.0;
 sq1_envAdd[328] = 0.0;
 sq1_envAdd[329] = 0.0;
 sq1_envAdd[330] = 0.0;
 sq1_envAdd[331] = 0.0;
 sq1_envAdd[332] = 0.0;
 sq1_envAdd[333] = 0.0;
 sq1_envAdd[334] = 0.0;
 sq1_envAdd[335] = 0.0;
 sq1_envAdd[336] = 0.0;
 sq1_envAdd[337] = 0.0;
 sq1_envAdd[338] = 0.0;
 sq1_envAdd[339] = 0.0;
 sq1_envAdd[340] = 0.0;
 sq1_envAdd[341] = 0.0;
 sq1_envAdd[342] = 0.0;
 sq1_envAdd[343] = 0.0;
 sq1_envAdd[344] = 0.0;
 sq1_envAdd[345] = 0.0;
 sq1_envAdd[346] = 0.0;
 sq1_envAdd[347] = 0.0;
 sq1_envAdd[348] = 0.0;
 sq1_envAdd[349] = 0.0;
 sq1_envAdd[350] = 0.0;
 sq1_envAdd[351] = 0.0;
 sq1_envAdd[352] = 0.0;
 sq1_envAdd[353] = 0.0;
 sq1_envAdd[354] = 0.0;
 sq1_envAdd[355] = 0.0;
 sq1_envAdd[356] = 0.0;
 sq1_envAdd[357] = 0.0;
 sq1_envAdd[358] = 0.0;
 sq1_envAdd[359] = 0.0;
 sq1_envAdd[360] = 0.0;
 sq1_envAdd[361] = 0.0;
 sq1_envAdd[362] = 0.0;
 sq1_envAdd[363] = 0.0;
 sq1_envAdd[364] = 0.0;
 sq1_envAdd[365] = 0.0;
 sq1_envAdd[366] = 0.0;
 sq1_envAdd[367] = 0.0;
 sq1_envAdd[368] = 0.0;
 sq1_envAdd[369] = 0.0;
 sq1_envAdd[370] = 0.0;
 sq1_envAdd[371] = 0.0;
 sq1_envAdd[372] = 0.0;
 sq1_envAdd[373] = 0.0;
 sq1_envAdd[374] = 0.0;
 sq1_envAdd[375] = 0.0;
 sq1_envAdd[376] = 0.0;
 sq1_envAdd[377] = 0.0;
 sq1_envAdd[378] = 0.0;
 sq1_period[0] = 4.0;
 sq1_period[1] = 4.0;
 sq1_period[2] = 4.0;
 sq1_period[3] = 4.0;
 sq1_period[4] = 4.0;
 sq1_period[5] = 4.0;
 sq1_period[6] = 4.0;
 sq1_period[7] = 4.0;
 sq1_period[8] = 4.0;
 sq1_period[9] = 4.0;
 sq1_period[10] = 4.0;
 sq1_period[11] = 4.0;
 sq1_period[12] = 4.0;
 sq1_period[13] = 4.0;
 sq1_period[14] = 4.0;
 sq1_period[15] = 4.0;
 sq1_period[16] = 4.0;
 sq1_period[17] = 4.0;
 sq1_period[18] = 4.0;
 sq1_period[19] = 4.0;
 sq1_period[20] = 4.0;
 sq1_period[21] = 4.0;
 sq1_period[22] = 4.0;
 sq1_period[23] = 4.0;
 sq1_period[24] = 4.0;
 sq1_period[25] = 4.0;
 sq1_period[26] = 4.0;
 sq1_period[27] = 4.0;
 sq1_period[28] = 4.0;
 sq1_period[29] = 4.0;
 sq1_period[30] = 4.0;
 sq1_period[31] = 4.0;
 sq1_period[32] = 4.0;
 sq1_period[33] = 4.0;
 sq1_period[34] = 4.0;
 sq1_period[35] = 4.0;
 sq1_period[36] = 4.0;
 sq1_period[37] = 4.0;
 sq1_period[38] = 4.0;
 sq1_period[39] = 4.0;
 sq1_period[40] = 4.0;
 sq1_period[41] = 4.0;
 sq1_period[42] = 4.0;
 sq1_period[43] = 4.0;
 sq1_period[44] = 4.0;
 sq1_period[45] = 4.0;
 sq1_period[46] = 4.0;
 sq1_period[47] = 4.0;
 sq1_period[48] = 4.0;
 sq1_period[49] = 4.0;
 sq1_period[50] = 4.0;
 sq1_period[51] = 4.0;
 sq1_period[52] = 4.0;
 sq1_period[53] = 4.0;
 sq1_period[54] = 4.0;
 sq1_period[55] = 4.0;
 sq1_period[56] = 4.0;
 sq1_period[57] = 4.0;
 sq1_period[58] = 4.0;
 sq1_period[59] = 4.0;
 sq1_period[60] = 4.0;
 sq1_period[61] = 4.0;
 sq1_period[62] = 4.0;
 sq1_period[63] = 4.0;
 sq1_period[64] = 4.0;
 sq1_period[65] = 4.0;
 sq1_period[66] = 4.0;
 sq1_period[67] = 4.0;
 sq1_period[68] = 4.0;
 sq1_period[69] = 4.0;
 sq1_period[70] = 4.0;
 sq1_period[71] = 4.0;
 sq1_period[72] = 4.0;
 sq1_period[73] = 4.0;
 sq1_period[74] = 4.0;
 sq1_period[75] = 4.0;
 sq1_period[76] = 4.0;
 sq1_period[77] = 4.0;
 sq1_period[78] = 4.0;
 sq1_period[79] = 4.0;
 sq1_period[80] = 4.0;
 sq1_period[81] = 4.0;
 sq1_period[82] = 4.0;
 sq1_period[83] = 4.0;
 sq1_period[84] = 4.0;
 sq1_period[85] = 4.0;
 sq1_period[86] = 4.0;
 sq1_period[87] = 4.0;
 sq1_period[88] = 4.0;
 sq1_period[89] = 4.0;
 sq1_period[90] = 4.0;
 sq1_period[91] = 4.0;
 sq1_period[92] = 4.0;
 sq1_period[93] = 4.0;
 sq1_period[94] = 4.0;
 sq1_period[95] = 4.0;
 sq1_period[96] = 4.0;
 sq1_period[97] = 4.0;
 sq1_period[98] = 4.0;
 sq1_period[99] = 4.0;
 sq1_period[100] = 4.0;
 sq1_period[101] = 4.0;
 sq1_period[102] = 4.0;
 sq1_period[103] = 4.0;
 sq1_period[104] = 4.0;
 sq1_period[105] = 4.0;
 sq1_period[106] = 4.0;
 sq1_period[107] = 4.0;
 sq1_period[108] = 4.0;
 sq1_period[109] = 4.0;
 sq1_period[110] = 4.0;
 sq1_period[111] = 4.0;
 sq1_period[112] = 4.0;
 sq1_period[113] = 4.0;
 sq1_period[114] = 4.0;
 sq1_period[115] = 4.0;
 sq1_period[116] = 4.0;
 sq1_period[117] = 4.0;
 sq1_period[118] = 4.0;
 sq1_period[119] = 4.0;
 sq1_period[120] = 4.0;
 sq1_period[121] = 4.0;
 sq1_period[122] = 4.0;
 sq1_period[123] = 4.0;
 sq1_period[124] = 4.0;
 sq1_period[125] = 4.0;
 sq1_period[126] = 4.0;
 sq1_period[127] = 4.0;
 sq1_period[128] = 4.0;
 sq1_period[129] = 4.0;
 sq1_period[130] = 4.0;
 sq1_period[131] = 4.0;
 sq1_period[132] = 4.0;
 sq1_period[133] = 4.0;
 sq1_period[134] = 4.0;
 sq1_period[135] = 4.0;
 sq1_period[136] = 4.0;
 sq1_period[137] = 4.0;
 sq1_period[138] = 4.0;
 sq1_period[139] = 4.0;
 sq1_period[140] = 4.0;
 sq1_period[141] = 4.0;
 sq1_period[142] = 4.0;
 sq1_period[143] = 4.0;
 sq1_period[144] = 4.0;
 sq1_period[145] = 4.0;
 sq1_period[146] = 4.0;
 sq1_period[147] = 4.0;
 sq1_period[148] = 4.0;
 sq1_period[149] = 4.0;
 sq1_period[150] = 4.0;
 sq1_period[151] = 4.0;
 sq1_period[152] = 4.0;
 sq1_period[153] = 4.0;
 sq1_period[154] = 4.0;
 sq1_period[155] = 4.0;
 sq1_period[156] = 4.0;
 sq1_period[157] = 4.0;
 sq1_period[158] = 4.0;
 sq1_period[159] = 4.0;
 sq1_period[160] = 4.0;
 sq1_period[161] = 4.0;
 sq1_period[162] = 4.0;
 sq1_period[163] = 4.0;
 sq1_period[164] = 4.0;
 sq1_period[165] = 4.0;
 sq1_period[166] = 4.0;
 sq1_period[167] = 4.0;
 sq1_period[168] = 4.0;
 sq1_period[169] = 4.0;
 sq1_period[170] = 4.0;
 sq1_period[171] = 4.0;
 sq1_period[172] = 4.0;
 sq1_period[173] = 4.0;
 sq1_period[174] = 4.0;
 sq1_period[175] = 4.0;
 sq1_period[176] = 4.0;
 sq1_period[177] = 4.0;
 sq1_period[178] = 4.0;
 sq1_period[179] = 4.0;
 sq1_period[180] = 4.0;
 sq1_period[181] = 4.0;
 sq1_period[182] = 4.0;
 sq1_period[183] = 4.0;
 sq1_period[184] = 4.0;
 sq1_period[185] = 4.0;
 sq1_period[186] = 4.0;
 sq1_period[187] = 4.0;
 sq1_period[188] = 4.0;
 sq1_period[189] = 4.0;
 sq1_period[190] = 4.0;
 sq1_period[191] = 4.0;
 sq1_period[192] = 4.0;
 sq1_period[193] = 4.0;
 sq1_period[194] = 4.0;
 sq1_period[195] = 4.0;
 sq1_period[196] = 4.0;
 sq1_period[197] = 4.0;
 sq1_period[198] = 4.0;
 sq1_period[199] = 4.0;
 sq1_period[200] = 4.0;
 sq1_period[201] = 4.0;
 sq1_period[202] = 4.0;
 sq1_period[203] = 4.0;
 sq1_period[204] = 4.0;
 sq1_period[205] = 4.0;
 sq1_period[206] = 4.0;
 sq1_period[207] = 4.0;
 sq1_period[208] = 4.0;
 sq1_period[209] = 4.0;
 sq1_period[210] = 4.0;
 sq1_period[211] = 4.0;
 sq1_period[212] = 4.0;
 sq1_period[213] = 4.0;
 sq1_period[214] = 4.0;
 sq1_period[215] = 4.0;
 sq1_period[216] = 4.0;
 sq1_period[217] = 4.0;
 sq1_period[218] = 4.0;
 sq1_period[219] = 4.0;
 sq1_period[220] = 4.0;
 sq1_period[221] = 4.0;
 sq1_period[222] = 4.0;
 sq1_period[223] = 4.0;
 sq1_period[224] = 4.0;
 sq1_period[225] = 4.0;
 sq1_period[226] = 4.0;
 sq1_period[227] = 4.0;
 sq1_period[228] = 4.0;
 sq1_period[229] = 4.0;
 sq1_period[230] = 4.0;
 sq1_period[231] = 4.0;
 sq1_period[232] = 4.0;
 sq1_period[233] = 4.0;
 sq1_period[234] = 4.0;
 sq1_period[235] = 4.0;
 sq1_period[236] = 4.0;
 sq1_period[237] = 4.0;
 sq1_period[238] = 4.0;
 sq1_period[239] = 4.0;
 sq1_period[240] = 4.0;
 sq1_period[241] = 4.0;
 sq1_period[242] = 4.0;
 sq1_period[243] = 4.0;
 sq1_period[244] = 4.0;
 sq1_period[245] = 4.0;
 sq1_period[246] = 4.0;
 sq1_period[247] = 4.0;
 sq1_period[248] = 4.0;
 sq1_period[249] = 4.0;
 sq1_period[250] = 4.0;
 sq1_period[251] = 4.0;
 sq1_period[252] = 4.0;
 sq1_period[253] = 4.0;
 sq1_period[254] = 4.0;
 sq1_period[255] = 4.0;
 sq1_period[256] = 4.0;
 sq1_period[257] = 4.0;
 sq1_period[258] = 4.0;
 sq1_period[259] = 4.0;
 sq1_period[260] = 4.0;
 sq1_period[261] = 4.0;
 sq1_period[262] = 4.0;
 sq1_period[263] = 4.0;
 sq1_period[264] = 4.0;
 sq1_period[265] = 4.0;
 sq1_period[266] = 4.0;
 sq1_period[267] = 4.0;
 sq1_period[268] = 4.0;
 sq1_period[269] = 4.0;
 sq1_period[270] = 4.0;
 sq1_period[271] = 4.0;
 sq1_period[272] = 4.0;
 sq1_period[273] = 4.0;
 sq1_period[274] = 4.0;
 sq1_period[275] = 4.0;
 sq1_period[276] = 4.0;
 sq1_period[277] = 4.0;
 sq1_period[278] = 4.0;
 sq1_period[279] = 4.0;
 sq1_period[280] = 4.0;
 sq1_period[281] = 4.0;
 sq1_period[282] = 4.0;
 sq1_period[283] = 4.0;
 sq1_period[284] = 4.0;
 sq1_period[285] = 4.0;
 sq1_period[286] = 4.0;
 sq1_period[287] = 4.0;
 sq1_period[288] = 4.0;
 sq1_period[289] = 4.0;
 sq1_period[290] = 4.0;
 sq1_period[291] = 4.0;
 sq1_period[292] = 4.0;
 sq1_period[293] = 4.0;
 sq1_period[294] = 4.0;
 sq1_period[295] = 4.0;
 sq1_period[296] = 4.0;
 sq1_period[297] = 4.0;
 sq1_period[298] = 4.0;
 sq1_period[299] = 4.0;
 sq1_period[300] = 4.0;
 sq1_period[301] = 4.0;
 sq1_period[302] = 4.0;
 sq1_period[303] = 4.0;
 sq1_period[304] = 4.0;
 sq1_period[305] = 4.0;
 sq1_period[306] = 4.0;
 sq1_period[307] = 4.0;
 sq1_period[308] = 4.0;
 sq1_period[309] = 4.0;
 sq1_period[310] = 4.0;
 sq1_period[311] = 4.0;
 sq1_period[312] = 4.0;
 sq1_period[313] = 4.0;
 sq1_period[314] = 4.0;
 sq1_period[315] = 4.0;
 sq1_period[316] = 4.0;
 sq1_period[317] = 4.0;
 sq1_period[318] = 4.0;
 sq1_period[319] = 4.0;
 sq1_period[320] = 4.0;
 sq1_period[321] = 4.0;
 sq1_period[322] = 4.0;
 sq1_period[323] = 4.0;
 sq1_period[324] = 4.0;
 sq1_period[325] = 4.0;
 sq1_period[326] = 4.0;
 sq1_period[327] = 4.0;
 sq1_period[328] = 4.0;
 sq1_period[329] = 4.0;
 sq1_period[330] = 4.0;
 sq1_period[331] = 4.0;
 sq1_period[332] = 4.0;
 sq1_period[333] = 4.0;
 sq1_period[334] = 4.0;
 sq1_period[335] = 4.0;
 sq1_period[336] = 4.0;
 sq1_period[337] = 4.0;
 sq1_period[338] = 4.0;
 sq1_period[339] = 4.0;
 sq1_period[340] = 4.0;
 sq1_period[341] = 4.0;
 sq1_period[342] = 4.0;
 sq1_period[343] = 4.0;
 sq1_period[344] = 4.0;
 sq1_period[345] = 4.0;
 sq1_period[346] = 4.0;
 sq1_period[347] = 4.0;
 sq1_period[348] = 4.0;
 sq1_period[349] = 4.0;
 sq1_period[350] = 4.0;
 sq1_period[351] = 4.0;
 sq1_period[352] = 4.0;
 sq1_period[353] = 4.0;
 sq1_period[354] = 4.0;
 sq1_period[355] = 4.0;
 sq1_period[356] = 4.0;
 sq1_period[357] = 4.0;
 sq1_period[358] = 4.0;
 sq1_period[359] = 4.0;
 sq1_period[360] = 4.0;
 sq1_period[361] = 4.0;
 sq1_period[362] = 4.0;
 sq1_period[363] = 4.0;
 sq1_period[364] = 4.0;
 sq1_period[365] = 4.0;
 sq1_period[366] = 4.0;
 sq1_period[367] = 4.0;
 sq1_period[368] = 4.0;
 sq1_period[369] = 4.0;
 sq1_period[370] = 4.0;
 sq1_period[371] = 4.0;
 sq1_period[372] = 4.0;
 sq1_period[373] = 4.0;
 sq1_period[374] = 4.0;
 sq1_period[375] = 4.0;
 sq1_period[376] = 4.0;
 sq1_period[377] = 4.0;
 sq1_period[378] = 4.0;
 sq1_freq[0] = 1714;
 sq1_freq[1] = 1714;
 sq1_freq[2] = 1714;
 sq1_freq[3] = 1714;
 sq1_freq[4] = 1714;
 sq1_freq[5] = 1714;
 sq1_freq[6] = 1714;
 sq1_freq[7] = 1714;
 sq1_freq[8] = 1714;
 sq1_freq[9] = 1714;
 sq1_freq[10] = 1714;
 sq1_freq[11] = 1714;
 sq1_freq[12] = 1602;
 sq1_freq[13] = 1602;
 sq1_freq[14] = 1602;
 sq1_freq[15] = 1602;
 sq1_freq[16] = 1602;
 sq1_freq[17] = 1602;
 sq1_freq[18] = 1602;
 sq1_freq[19] = 1602;
 sq1_freq[20] = 1602;
 sq1_freq[21] = 1602;
 sq1_freq[22] = 1602;
 sq1_freq[23] = 1602;
 sq1_freq[24] = 1602;
 sq1_freq[25] = 1602;
 sq1_freq[26] = 1602;
 sq1_freq[27] = 1602;
 sq1_freq[28] = 1602;
 sq1_freq[29] = 1602;
 sq1_freq[30] = 1714;
 sq1_freq[31] = 1714;
 sq1_freq[32] = 1714;
 sq1_freq[33] = 1714;
 sq1_freq[34] = 1714;
 sq1_freq[35] = 1714;
 sq1_freq[36] = 1714;
 sq1_freq[37] = 1714;
 sq1_freq[38] = 1714;
 sq1_freq[39] = 1750;
 sq1_freq[40] = 1750;
 sq1_freq[41] = 1750;
 sq1_freq[42] = 1783;
 sq1_freq[43] = 1783;
 sq1_freq[44] = 1783;
 sq1_freq[45] = 1798;
 sq1_freq[46] = 1798;
 sq1_freq[47] = 1798;
 sq1_freq[48] = 1825;
 sq1_freq[49] = 1825;
 sq1_freq[50] = 1825;
 sq1_freq[51] = 1825;
 sq1_freq[52] = 1825;
 sq1_freq[53] = 1825;
 sq1_freq[54] = 1825;
 sq1_freq[55] = 1825;
 sq1_freq[56] = 1825;
 sq1_freq[57] = 1825;
 sq1_freq[58] = 1825;
 sq1_freq[59] = 1825;
 sq1_freq[60] = 1825;
 sq1_freq[61] = 1825;
 sq1_freq[62] = 1825;
 sq1_freq[63] = 1825;
 sq1_freq[64] = 1825;
 sq1_freq[65] = 1825;
 sq1_freq[66] = 1825;
 sq1_freq[67] = 1825;
 sq1_freq[68] = 1825;
 sq1_freq[69] = 1825;
 sq1_freq[70] = 1825;
 sq1_freq[71] = 1825;
 sq1_freq[72] = 1825;
 sq1_freq[73] = 1825;
 sq1_freq[74] = 1825;
 sq1_freq[75] = 1825;
 sq1_freq[76] = 1825;
 sq1_freq[77] = 1825;
 sq1_freq[78] = 1825;
 sq1_freq[79] = 1825;
 sq1_freq[80] = 1825;
 sq1_freq[81] = 1825;
 sq1_freq[82] = 1825;
 sq1_freq[83] = 1825;
 sq1_freq[84] = 1825;
 sq1_freq[85] = 1825;
 sq1_freq[86] = 1825;
 sq1_freq[87] = 1825;
 sq1_freq[88] = 1837;
 sq1_freq[89] = 1837;
 sq1_freq[90] = 1837;
 sq1_freq[91] = 1837;
 sq1_freq[92] = 1860;
 sq1_freq[93] = 1860;
 sq1_freq[94] = 1860;
 sq1_freq[95] = 1860;
 sq1_freq[96] = 1881;
 sq1_freq[97] = 1881;
 sq1_freq[98] = 1881;
 sq1_freq[99] = 1881;
 sq1_freq[100] = 1881;
 sq1_freq[101] = 1881;
 sq1_freq[102] = 1881;
 sq1_freq[103] = 1881;
 sq1_freq[104] = 1881;
 sq1_freq[105] = 1881;
 sq1_freq[106] = 1881;
 sq1_freq[107] = 1881;
 sq1_freq[108] = 1881;
 sq1_freq[109] = 1881;
 sq1_freq[110] = 1881;
 sq1_freq[111] = 1881;
 sq1_freq[112] = 1881;
 sq1_freq[113] = 1881;
 sq1_freq[114] = 1881;
 sq1_freq[115] = 1881;
 sq1_freq[116] = 1881;
 sq1_freq[117] = 1881;
 sq1_freq[118] = 1881;
 sq1_freq[119] = 1881;
 sq1_freq[120] = 1881;
 sq1_freq[121] = 1881;
 sq1_freq[122] = 1881;
 sq1_freq[123] = 1881;
 sq1_freq[124] = 1881;
 sq1_freq[125] = 1881;
 sq1_freq[126] = 1881;
 sq1_freq[127] = 1881;
 sq1_freq[128] = 1881;
 sq1_freq[129] = 1881;
 sq1_freq[130] = 1881;
 sq1_freq[131] = 1881;
 sq1_freq[132] = 1881;
 sq1_freq[133] = 1881;
 sq1_freq[134] = 1881;
 sq1_freq[135] = 1881;
 sq1_freq[136] = 1860;
 sq1_freq[137] = 1860;
 sq1_freq[138] = 1860;
 sq1_freq[139] = 1860;
 sq1_freq[140] = 1837;
 sq1_freq[141] = 1837;
 sq1_freq[142] = 1837;
 sq1_freq[143] = 1837;
 sq1_freq[144] = 1860;
 sq1_freq[145] = 1860;
 sq1_freq[146] = 1860;
 sq1_freq[147] = 1860;
 sq1_freq[148] = 1860;
 sq1_freq[149] = 1860;
 sq1_freq[150] = 1860;
 sq1_freq[151] = 1860;
 sq1_freq[152] = 1837;
 sq1_freq[153] = 1837;
 sq1_freq[154] = 1837;
 sq1_freq[155] = 1837;
 sq1_freq[156] = 1825;
 sq1_freq[157] = 1825;
 sq1_freq[158] = 1825;
 sq1_freq[159] = 1825;
 sq1_freq[160] = 1825;
 sq1_freq[161] = 1825;
 sq1_freq[162] = 1825;
 sq1_freq[163] = 1825;
 sq1_freq[164] = 1825;
 sq1_freq[165] = 1825;
 sq1_freq[166] = 1825;
 sq1_freq[167] = 1825;
 sq1_freq[168] = 1825;
 sq1_freq[169] = 1825;
 sq1_freq[170] = 1825;
 sq1_freq[171] = 1825;
 sq1_freq[172] = 1825;
 sq1_freq[173] = 1825;
 sq1_freq[174] = 1825;
 sq1_freq[175] = 1825;
 sq1_freq[176] = 1825;
 sq1_freq[177] = 1825;
 sq1_freq[178] = 1825;
 sq1_freq[179] = 1825;
 sq1_freq[180] = 1825;
 sq1_freq[181] = 1825;
 sq1_freq[182] = 1825;
 sq1_freq[183] = 1825;
 sq1_freq[184] = 1825;
 sq1_freq[185] = 1825;
 sq1_freq[186] = 1825;
 sq1_freq[187] = 1825;
 sq1_freq[188] = 1825;
 sq1_freq[189] = 1825;
 sq1_freq[190] = 1825;
 sq1_freq[191] = 1825;
 sq1_freq[192] = 1798;
 sq1_freq[193] = 1798;
 sq1_freq[194] = 1798;
 sq1_freq[195] = 1798;
 sq1_freq[196] = 1798;
 sq1_freq[197] = 1798;
 sq1_freq[198] = 1798;
 sq1_freq[199] = 1798;
 sq1_freq[200] = 1798;
 sq1_freq[201] = 1825;
 sq1_freq[202] = 1825;
 sq1_freq[203] = 1825;
 sq1_freq[204] = 1837;
 sq1_freq[205] = 1837;
 sq1_freq[206] = 1837;
 sq1_freq[207] = 1837;
 sq1_freq[208] = 1837;
 sq1_freq[209] = 1837;
 sq1_freq[210] = 1837;
 sq1_freq[211] = 1837;
 sq1_freq[212] = 1837;
 sq1_freq[213] = 1837;
 sq1_freq[214] = 1837;
 sq1_freq[215] = 1837;
 sq1_freq[216] = 1837;
 sq1_freq[217] = 1837;
 sq1_freq[218] = 1837;
 sq1_freq[219] = 1837;
 sq1_freq[220] = 1837;
 sq1_freq[221] = 1837;
 sq1_freq[222] = 1837;
 sq1_freq[223] = 1837;
 sq1_freq[224] = 1837;
 sq1_freq[225] = 1837;
 sq1_freq[226] = 1837;
 sq1_freq[227] = 1837;
 sq1_freq[228] = 1825;
 sq1_freq[229] = 1825;
 sq1_freq[230] = 1825;
 sq1_freq[231] = 1825;
 sq1_freq[232] = 1825;
 sq1_freq[233] = 1825;
 sq1_freq[234] = 1798;
 sq1_freq[235] = 1798;
 sq1_freq[236] = 1798;
 sq1_freq[237] = 1798;
 sq1_freq[238] = 1798;
 sq1_freq[239] = 1798;
 sq1_freq[240] = 1767;
 sq1_freq[241] = 1767;
 sq1_freq[242] = 1767;
 sq1_freq[243] = 1767;
 sq1_freq[244] = 1767;
 sq1_freq[245] = 1767;
 sq1_freq[246] = 1767;
 sq1_freq[247] = 1767;
 sq1_freq[248] = 1767;
 sq1_freq[249] = 1798;
 sq1_freq[250] = 1798;
 sq1_freq[251] = 1798;
 sq1_freq[252] = 1825;
 sq1_freq[253] = 1825;
 sq1_freq[254] = 1825;
 sq1_freq[255] = 1825;
 sq1_freq[256] = 1825;
 sq1_freq[257] = 1825;
 sq1_freq[258] = 1825;
 sq1_freq[259] = 1825;
 sq1_freq[260] = 1825;
 sq1_freq[261] = 1825;
 sq1_freq[262] = 1825;
 sq1_freq[263] = 1825;
 sq1_freq[264] = 1825;
 sq1_freq[265] = 1825;
 sq1_freq[266] = 1825;
 sq1_freq[267] = 1825;
 sq1_freq[268] = 1825;
 sq1_freq[269] = 1825;
 sq1_freq[270] = 1825;
 sq1_freq[271] = 1825;
 sq1_freq[272] = 1825;
 sq1_freq[273] = 1825;
 sq1_freq[274] = 1825;
 sq1_freq[275] = 1825;
 sq1_freq[276] = 1798;
 sq1_freq[277] = 1798;
 sq1_freq[278] = 1798;
 sq1_freq[279] = 1798;
 sq1_freq[280] = 1798;
 sq1_freq[281] = 1798;
 sq1_freq[282] = 1767;
 sq1_freq[283] = 1767;
 sq1_freq[284] = 1767;
 sq1_freq[285] = 1767;
 sq1_freq[286] = 1767;
 sq1_freq[287] = 1767;
 sq1_freq[288] = 1750;
 sq1_freq[289] = 1750;
 sq1_freq[290] = 1750;
 sq1_freq[291] = 1750;
 sq1_freq[292] = 1750;
 sq1_freq[293] = 1750;
 sq1_freq[294] = 1750;
 sq1_freq[295] = 1750;
 sq1_freq[296] = 1750;
 sq1_freq[297] = 1783;
 sq1_freq[298] = 1783;
 sq1_freq[299] = 1783;
 sq1_freq[300] = 1812;
 sq1_freq[301] = 1812;
 sq1_freq[302] = 1812;
 sq1_freq[303] = 1812;
 sq1_freq[304] = 1812;
 sq1_freq[305] = 1812;
 sq1_freq[306] = 1812;
 sq1_freq[307] = 1812;
 sq1_freq[308] = 1812;
 sq1_freq[309] = 1812;
 sq1_freq[310] = 1812;
 sq1_freq[311] = 1812;
 sq1_freq[312] = 1812;
 sq1_freq[313] = 1812;
 sq1_freq[314] = 1812;
 sq1_freq[315] = 1812;
 sq1_freq[316] = 1812;
 sq1_freq[317] = 1812;
 sq1_freq[318] = 1812;
 sq1_freq[319] = 1812;
 sq1_freq[320] = 1812;
 sq1_freq[321] = 1812;
 sq1_freq[322] = 1812;
 sq1_freq[323] = 1812;
 sq1_freq[324] = 1849;
 sq1_freq[325] = 1849;
 sq1_freq[326] = 1849;
 sq1_freq[327] = 1849;
 sq1_freq[328] = 1849;
 sq1_freq[329] = 1849;
 sq1_freq[330] = 1849;
 sq1_freq[331] = 1849;
 sq1_freq[332] = 1849;
 sq1_freq[333] = 1849;
 sq1_freq[334] = 1849;
 sq1_freq[335] = 1849;
 sq1_freq[336] = 1825;
 sq1_freq[337] = 1825;
 sq1_freq[338] = 1825;
 sq1_freq[339] = 1825;
 sq1_freq[340] = 1825;
 sq1_freq[341] = 1825;
 sq1_freq[342] = 1825;
 sq1_freq[343] = 1825;
 sq1_freq[344] = 1825;
 sq1_freq[345] = 1825;
 sq1_freq[346] = 1825;
 sq1_freq[347] = 1825;
 sq1_freq[348] = 1825;
 sq1_freq[349] = 1825;
 sq1_freq[350] = 1825;
 sq1_freq[351] = 1825;
 sq1_freq[352] = 1825;
 sq1_freq[353] = 1825;
 sq1_freq[354] = 1825;
 sq1_freq[355] = 1825;
 sq1_freq[356] = 1825;
 sq1_freq[357] = 1825;
 sq1_freq[358] = 1825;
 sq1_freq[359] = 1825;
 sq1_freq[360] = 1825;
 sq1_freq[361] = 1825;
 sq1_freq[362] = 1825;
 sq1_freq[363] = 1825;
 sq1_freq[364] = 1825;
 sq1_freq[365] = 1825;
 sq1_freq[366] = 1825;
 sq1_freq[367] = 1825;
 sq1_freq[368] = 1825;
 sq1_freq[369] = 1825;
 sq1_freq[370] = 1825;
 sq1_freq[371] = 1825;
 sq1_freq[372] = 1825;
 sq1_freq[373] = 1825;
 sq1_freq[374] = 1825;
 sq1_freq[375] = 1825;
 sq1_freq[376] = 1825;
 sq1_freq[377] = 1825;
 sq1_freq[378] = 1825;
 sq1_trigger[0] = 1.0;
 sq1_trigger[1] = 0;
 sq1_trigger[2] = 0;
 sq1_trigger[3] = 0;
 sq1_trigger[4] = 0;
 sq1_trigger[5] = 0;
 sq1_trigger[6] = 0;
 sq1_trigger[7] = 0;
 sq1_trigger[8] = 0;
 sq1_trigger[9] = 0;
 sq1_trigger[10] = 0;
 sq1_trigger[11] = 0;
 sq1_trigger[12] = 1.0;
 sq1_trigger[13] = 0;
 sq1_trigger[14] = 0;
 sq1_trigger[15] = 0;
 sq1_trigger[16] = 0;
 sq1_trigger[17] = 0;
 sq1_trigger[18] = 0;
 sq1_trigger[19] = 0;
 sq1_trigger[20] = 0;
 sq1_trigger[21] = 0;
 sq1_trigger[22] = 0;
 sq1_trigger[23] = 0;
 sq1_trigger[24] = 0;
 sq1_trigger[25] = 0;
 sq1_trigger[26] = 0;
 sq1_trigger[27] = 0;
 sq1_trigger[28] = 0;
 sq1_trigger[29] = 0;
 sq1_trigger[30] = 1.0;
 sq1_trigger[31] = 0;
 sq1_trigger[32] = 0;
 sq1_trigger[33] = 0;
 sq1_trigger[34] = 0;
 sq1_trigger[35] = 0;
 sq1_trigger[36] = 1.0;
 sq1_trigger[37] = 0;
 sq1_trigger[38] = 0;
 sq1_trigger[39] = 1.0;
 sq1_trigger[40] = 0;
 sq1_trigger[41] = 0;
 sq1_trigger[42] = 1.0;
 sq1_trigger[43] = 0;
 sq1_trigger[44] = 0;
 sq1_trigger[45] = 1.0;
 sq1_trigger[46] = 0;
 sq1_trigger[47] = 0;
 sq1_trigger[48] = 1.0;
 sq1_trigger[49] = 0;
 sq1_trigger[50] = 0;
 sq1_trigger[51] = 0;
 sq1_trigger[52] = 0;
 sq1_trigger[53] = 0;
 sq1_trigger[54] = 0;
 sq1_trigger[55] = 0;
 sq1_trigger[56] = 0;
 sq1_trigger[57] = 0;
 sq1_trigger[58] = 0;
 sq1_trigger[59] = 0;
 sq1_trigger[60] = 0;
 sq1_trigger[61] = 0;
 sq1_trigger[62] = 0;
 sq1_trigger[63] = 0;
 sq1_trigger[64] = 0;
 sq1_trigger[65] = 0;
 sq1_trigger[66] = 0;
 sq1_trigger[67] = 0;
 sq1_trigger[68] = 0;
 sq1_trigger[69] = 0;
 sq1_trigger[70] = 0;
 sq1_trigger[71] = 0;
 sq1_trigger[72] = 0;
 sq1_trigger[73] = 0;
 sq1_trigger[74] = 0;
 sq1_trigger[75] = 0;
 sq1_trigger[76] = 0;
 sq1_trigger[77] = 0;
 sq1_trigger[78] = 1.0;
 sq1_trigger[79] = 0;
 sq1_trigger[80] = 0;
 sq1_trigger[81] = 0;
 sq1_trigger[82] = 0;
 sq1_trigger[83] = 0;
 sq1_trigger[84] = 1.0;
 sq1_trigger[85] = 0;
 sq1_trigger[86] = 0;
 sq1_trigger[87] = 0;
 sq1_trigger[88] = 1.0;
 sq1_trigger[89] = 0;
 sq1_trigger[90] = 0;
 sq1_trigger[91] = 0;
 sq1_trigger[92] = 1.0;
 sq1_trigger[93] = 0;
 sq1_trigger[94] = 0;
 sq1_trigger[95] = 0;
 sq1_trigger[96] = 1.0;
 sq1_trigger[97] = 0;
 sq1_trigger[98] = 0;
 sq1_trigger[99] = 0;
 sq1_trigger[100] = 0;
 sq1_trigger[101] = 0;
 sq1_trigger[102] = 0;
 sq1_trigger[103] = 0;
 sq1_trigger[104] = 0;
 sq1_trigger[105] = 0;
 sq1_trigger[106] = 0;
 sq1_trigger[107] = 0;
 sq1_trigger[108] = 0;
 sq1_trigger[109] = 0;
 sq1_trigger[110] = 0;
 sq1_trigger[111] = 0;
 sq1_trigger[112] = 0;
 sq1_trigger[113] = 0;
 sq1_trigger[114] = 0;
 sq1_trigger[115] = 0;
 sq1_trigger[116] = 0;
 sq1_trigger[117] = 0;
 sq1_trigger[118] = 0;
 sq1_trigger[119] = 0;
 sq1_trigger[120] = 0;
 sq1_trigger[121] = 0;
 sq1_trigger[122] = 0;
 sq1_trigger[123] = 0;
 sq1_trigger[124] = 1.0;
 sq1_trigger[125] = 0;
 sq1_trigger[126] = 0;
 sq1_trigger[127] = 0;
 sq1_trigger[128] = 1.0;
 sq1_trigger[129] = 0;
 sq1_trigger[130] = 0;
 sq1_trigger[131] = 0;
 sq1_trigger[132] = 1.0;
 sq1_trigger[133] = 0;
 sq1_trigger[134] = 0;
 sq1_trigger[135] = 0;
 sq1_trigger[136] = 1.0;
 sq1_trigger[137] = 0;
 sq1_trigger[138] = 0;
 sq1_trigger[139] = 0;
 sq1_trigger[140] = 1.0;
 sq1_trigger[141] = 0;
 sq1_trigger[142] = 0;
 sq1_trigger[143] = 0;
 sq1_trigger[144] = 1.0;
 sq1_trigger[145] = 0;
 sq1_trigger[146] = 0;
 sq1_trigger[147] = 0;
 sq1_trigger[148] = 0;
 sq1_trigger[149] = 0;
 sq1_trigger[150] = 0;
 sq1_trigger[151] = 0;
 sq1_trigger[152] = 1.0;
 sq1_trigger[153] = 0;
 sq1_trigger[154] = 0;
 sq1_trigger[155] = 0;
 sq1_trigger[156] = 1.0;
 sq1_trigger[157] = 0;
 sq1_trigger[158] = 0;
 sq1_trigger[159] = 0;
 sq1_trigger[160] = 0;
 sq1_trigger[161] = 0;
 sq1_trigger[162] = 0;
 sq1_trigger[163] = 0;
 sq1_trigger[164] = 0;
 sq1_trigger[165] = 0;
 sq1_trigger[166] = 0;
 sq1_trigger[167] = 0;
 sq1_trigger[168] = 0;
 sq1_trigger[169] = 0;
 sq1_trigger[170] = 0;
 sq1_trigger[171] = 0;
 sq1_trigger[172] = 0;
 sq1_trigger[173] = 0;
 sq1_trigger[174] = 0;
 sq1_trigger[175] = 0;
 sq1_trigger[176] = 0;
 sq1_trigger[177] = 0;
 sq1_trigger[178] = 0;
 sq1_trigger[179] = 0;
 sq1_trigger[180] = 1.0;
 sq1_trigger[181] = 0;
 sq1_trigger[182] = 0;
 sq1_trigger[183] = 0;
 sq1_trigger[184] = 0;
 sq1_trigger[185] = 0;
 sq1_trigger[186] = 0;
 sq1_trigger[187] = 0;
 sq1_trigger[188] = 0;
 sq1_trigger[189] = 0;
 sq1_trigger[190] = 0;
 sq1_trigger[191] = 0;
 sq1_trigger[192] = 1.0;
 sq1_trigger[193] = 0;
 sq1_trigger[194] = 0;
 sq1_trigger[195] = 0;
 sq1_trigger[196] = 0;
 sq1_trigger[197] = 0;
 sq1_trigger[198] = 1.0;
 sq1_trigger[199] = 0;
 sq1_trigger[200] = 0;
 sq1_trigger[201] = 1.0;
 sq1_trigger[202] = 0;
 sq1_trigger[203] = 0;
 sq1_trigger[204] = 1.0;
 sq1_trigger[205] = 0;
 sq1_trigger[206] = 0;
 sq1_trigger[207] = 0;
 sq1_trigger[208] = 0;
 sq1_trigger[209] = 0;
 sq1_trigger[210] = 0;
 sq1_trigger[211] = 0;
 sq1_trigger[212] = 0;
 sq1_trigger[213] = 0;
 sq1_trigger[214] = 0;
 sq1_trigger[215] = 0;
 sq1_trigger[216] = 0;
 sq1_trigger[217] = 0;
 sq1_trigger[218] = 0;
 sq1_trigger[219] = 0;
 sq1_trigger[220] = 0;
 sq1_trigger[221] = 0;
 sq1_trigger[222] = 0;
 sq1_trigger[223] = 0;
 sq1_trigger[224] = 0;
 sq1_trigger[225] = 0;
 sq1_trigger[226] = 0;
 sq1_trigger[227] = 0;
 sq1_trigger[228] = 1.0;
 sq1_trigger[229] = 0;
 sq1_trigger[230] = 0;
 sq1_trigger[231] = 0;
 sq1_trigger[232] = 0;
 sq1_trigger[233] = 0;
 sq1_trigger[234] = 1.0;
 sq1_trigger[235] = 0;
 sq1_trigger[236] = 0;
 sq1_trigger[237] = 0;
 sq1_trigger[238] = 0;
 sq1_trigger[239] = 0;
 sq1_trigger[240] = 1.0;
 sq1_trigger[241] = 0;
 sq1_trigger[242] = 0;
 sq1_trigger[243] = 0;
 sq1_trigger[244] = 0;
 sq1_trigger[245] = 0;
 sq1_trigger[246] = 1.0;
 sq1_trigger[247] = 0;
 sq1_trigger[248] = 0;
 sq1_trigger[249] = 1.0;
 sq1_trigger[250] = 0;
 sq1_trigger[251] = 0;
 sq1_trigger[252] = 1.0;
 sq1_trigger[253] = 0;
 sq1_trigger[254] = 0;
 sq1_trigger[255] = 0;
 sq1_trigger[256] = 0;
 sq1_trigger[257] = 0;
 sq1_trigger[258] = 0;
 sq1_trigger[259] = 0;
 sq1_trigger[260] = 0;
 sq1_trigger[261] = 0;
 sq1_trigger[262] = 0;
 sq1_trigger[263] = 0;
 sq1_trigger[264] = 0;
 sq1_trigger[265] = 0;
 sq1_trigger[266] = 0;
 sq1_trigger[267] = 0;
 sq1_trigger[268] = 0;
 sq1_trigger[269] = 0;
 sq1_trigger[270] = 0;
 sq1_trigger[271] = 0;
 sq1_trigger[272] = 0;
 sq1_trigger[273] = 0;
 sq1_trigger[274] = 0;
 sq1_trigger[275] = 0;
 sq1_trigger[276] = 1.0;
 sq1_trigger[277] = 0;
 sq1_trigger[278] = 0;
 sq1_trigger[279] = 0;
 sq1_trigger[280] = 0;
 sq1_trigger[281] = 0;
 sq1_trigger[282] = 1.0;
 sq1_trigger[283] = 0;
 sq1_trigger[284] = 0;
 sq1_trigger[285] = 0;
 sq1_trigger[286] = 0;
 sq1_trigger[287] = 0;
 sq1_trigger[288] = 1.0;
 sq1_trigger[289] = 0;
 sq1_trigger[290] = 0;
 sq1_trigger[291] = 0;
 sq1_trigger[292] = 0;
 sq1_trigger[293] = 0;
 sq1_trigger[294] = 1.0;
 sq1_trigger[295] = 0;
 sq1_trigger[296] = 0;
 sq1_trigger[297] = 1.0;
 sq1_trigger[298] = 0;
 sq1_trigger[299] = 0;
 sq1_trigger[300] = 1.0;
 sq1_trigger[301] = 0;
 sq1_trigger[302] = 0;
 sq1_trigger[303] = 0;
 sq1_trigger[304] = 0;
 sq1_trigger[305] = 0;
 sq1_trigger[306] = 0;
 sq1_trigger[307] = 0;
 sq1_trigger[308] = 0;
 sq1_trigger[309] = 0;
 sq1_trigger[310] = 0;
 sq1_trigger[311] = 0;
 sq1_trigger[312] = 0;
 sq1_trigger[313] = 0;
 sq1_trigger[314] = 0;
 sq1_trigger[315] = 0;
 sq1_trigger[316] = 0;
 sq1_trigger[317] = 0;
 sq1_trigger[318] = 0;
 sq1_trigger[319] = 0;
 sq1_trigger[320] = 0;
 sq1_trigger[321] = 0;
 sq1_trigger[322] = 0;
 sq1_trigger[323] = 0;
 sq1_trigger[324] = 1.0;
 sq1_trigger[325] = 0;
 sq1_trigger[326] = 0;
 sq1_trigger[327] = 0;
 sq1_trigger[328] = 0;
 sq1_trigger[329] = 0;
 sq1_trigger[330] = 0;
 sq1_trigger[331] = 0;
 sq1_trigger[332] = 0;
 sq1_trigger[333] = 0;
 sq1_trigger[334] = 0;
 sq1_trigger[335] = 0;
 sq1_trigger[336] = 1.0;
 sq1_trigger[337] = 0;
 sq1_trigger[338] = 0;
 sq1_trigger[339] = 0;
 sq1_trigger[340] = 0;
 sq1_trigger[341] = 0;
 sq1_trigger[342] = 0;
 sq1_trigger[343] = 0;
 sq1_trigger[344] = 0;
 sq1_trigger[345] = 0;
 sq1_trigger[346] = 0;
 sq1_trigger[347] = 0;
 sq1_trigger[348] = 0;
 sq1_trigger[349] = 0;
 sq1_trigger[350] = 0;
 sq1_trigger[351] = 0;
 sq1_trigger[352] = 0;
 sq1_trigger[353] = 0;
 sq1_trigger[354] = 0;
 sq1_trigger[355] = 0;
 sq1_trigger[356] = 0;
 sq1_trigger[357] = 0;
 sq1_trigger[358] = 0;
 sq1_trigger[359] = 0;
 sq1_trigger[360] = 0;
 sq1_trigger[361] = 0;
 sq1_trigger[362] = 0;
 sq1_trigger[363] = 0;
 sq1_trigger[364] = 0;
 sq1_trigger[365] = 0;
 sq1_trigger[366] = 0;
 sq1_trigger[367] = 0;
 sq1_trigger[368] = 0;
 sq1_trigger[369] = 0;
 sq1_trigger[370] = 0;
 sq1_trigger[371] = 0;
 sq1_trigger[372] = 0;
 sq1_trigger[373] = 0;
 sq1_trigger[374] = 0;
 sq1_trigger[375] = 0;
 sq1_trigger[376] = 0;
 sq1_trigger[377] = 0;
 sq1_trigger[378] = 0;
 sq1_lenEnable[0] = 1.0;
 sq1_lenEnable[1] = 1.0;
 sq1_lenEnable[2] = 1.0;
 sq1_lenEnable[3] = 1.0;
 sq1_lenEnable[4] = 1.0;
 sq1_lenEnable[5] = 1.0;
 sq1_lenEnable[6] = 1.0;
 sq1_lenEnable[7] = 1.0;
 sq1_lenEnable[8] = 1.0;
 sq1_lenEnable[9] = 1.0;
 sq1_lenEnable[10] = 1.0;
 sq1_lenEnable[11] = 1.0;
 sq1_lenEnable[12] = 1.0;
 sq1_lenEnable[13] = 1.0;
 sq1_lenEnable[14] = 1.0;
 sq1_lenEnable[15] = 1.0;
 sq1_lenEnable[16] = 1.0;
 sq1_lenEnable[17] = 1.0;
 sq1_lenEnable[18] = 1.0;
 sq1_lenEnable[19] = 1.0;
 sq1_lenEnable[20] = 1.0;
 sq1_lenEnable[21] = 1.0;
 sq1_lenEnable[22] = 1.0;
 sq1_lenEnable[23] = 1.0;
 sq1_lenEnable[24] = 1.0;
 sq1_lenEnable[25] = 1.0;
 sq1_lenEnable[26] = 1.0;
 sq1_lenEnable[27] = 1.0;
 sq1_lenEnable[28] = 1.0;
 sq1_lenEnable[29] = 1.0;
 sq1_lenEnable[30] = 1.0;
 sq1_lenEnable[31] = 1.0;
 sq1_lenEnable[32] = 1.0;
 sq1_lenEnable[33] = 1.0;
 sq1_lenEnable[34] = 1.0;
 sq1_lenEnable[35] = 1.0;
 sq1_lenEnable[36] = 1.0;
 sq1_lenEnable[37] = 1.0;
 sq1_lenEnable[38] = 1.0;
 sq1_lenEnable[39] = 1.0;
 sq1_lenEnable[40] = 1.0;
 sq1_lenEnable[41] = 1.0;
 sq1_lenEnable[42] = 1.0;
 sq1_lenEnable[43] = 1.0;
 sq1_lenEnable[44] = 1.0;
 sq1_lenEnable[45] = 1.0;
 sq1_lenEnable[46] = 1.0;
 sq1_lenEnable[47] = 1.0;
 sq1_lenEnable[48] = 1.0;
 sq1_lenEnable[49] = 1.0;
 sq1_lenEnable[50] = 1.0;
 sq1_lenEnable[51] = 1.0;
 sq1_lenEnable[52] = 1.0;
 sq1_lenEnable[53] = 1.0;
 sq1_lenEnable[54] = 1.0;
 sq1_lenEnable[55] = 1.0;
 sq1_lenEnable[56] = 1.0;
 sq1_lenEnable[57] = 1.0;
 sq1_lenEnable[58] = 1.0;
 sq1_lenEnable[59] = 1.0;
 sq1_lenEnable[60] = 1.0;
 sq1_lenEnable[61] = 1.0;
 sq1_lenEnable[62] = 1.0;
 sq1_lenEnable[63] = 1.0;
 sq1_lenEnable[64] = 1.0;
 sq1_lenEnable[65] = 1.0;
 sq1_lenEnable[66] = 1.0;
 sq1_lenEnable[67] = 1.0;
 sq1_lenEnable[68] = 1.0;
 sq1_lenEnable[69] = 1.0;
 sq1_lenEnable[70] = 1.0;
 sq1_lenEnable[71] = 1.0;
 sq1_lenEnable[72] = 1.0;
 sq1_lenEnable[73] = 1.0;
 sq1_lenEnable[74] = 1.0;
 sq1_lenEnable[75] = 1.0;
 sq1_lenEnable[76] = 1.0;
 sq1_lenEnable[77] = 1.0;
 sq1_lenEnable[78] = 1.0;
 sq1_lenEnable[79] = 1.0;
 sq1_lenEnable[80] = 1.0;
 sq1_lenEnable[81] = 1.0;
 sq1_lenEnable[82] = 1.0;
 sq1_lenEnable[83] = 1.0;
 sq1_lenEnable[84] = 1.0;
 sq1_lenEnable[85] = 1.0;
 sq1_lenEnable[86] = 1.0;
 sq1_lenEnable[87] = 1.0;
 sq1_lenEnable[88] = 1.0;
 sq1_lenEnable[89] = 1.0;
 sq1_lenEnable[90] = 1.0;
 sq1_lenEnable[91] = 1.0;
 sq1_lenEnable[92] = 1.0;
 sq1_lenEnable[93] = 1.0;
 sq1_lenEnable[94] = 1.0;
 sq1_lenEnable[95] = 1.0;
 sq1_lenEnable[96] = 1.0;
 sq1_lenEnable[97] = 1.0;
 sq1_lenEnable[98] = 1.0;
 sq1_lenEnable[99] = 1.0;
 sq1_lenEnable[100] = 1.0;
 sq1_lenEnable[101] = 1.0;
 sq1_lenEnable[102] = 1.0;
 sq1_lenEnable[103] = 1.0;
 sq1_lenEnable[104] = 1.0;
 sq1_lenEnable[105] = 1.0;
 sq1_lenEnable[106] = 1.0;
 sq1_lenEnable[107] = 1.0;
 sq1_lenEnable[108] = 1.0;
 sq1_lenEnable[109] = 1.0;
 sq1_lenEnable[110] = 1.0;
 sq1_lenEnable[111] = 1.0;
 sq1_lenEnable[112] = 1.0;
 sq1_lenEnable[113] = 1.0;
 sq1_lenEnable[114] = 1.0;
 sq1_lenEnable[115] = 1.0;
 sq1_lenEnable[116] = 1.0;
 sq1_lenEnable[117] = 1.0;
 sq1_lenEnable[118] = 1.0;
 sq1_lenEnable[119] = 1.0;
 sq1_lenEnable[120] = 1.0;
 sq1_lenEnable[121] = 1.0;
 sq1_lenEnable[122] = 1.0;
 sq1_lenEnable[123] = 1.0;
 sq1_lenEnable[124] = 1.0;
 sq1_lenEnable[125] = 1.0;
 sq1_lenEnable[126] = 1.0;
 sq1_lenEnable[127] = 1.0;
 sq1_lenEnable[128] = 1.0;
 sq1_lenEnable[129] = 1.0;
 sq1_lenEnable[130] = 1.0;
 sq1_lenEnable[131] = 1.0;
 sq1_lenEnable[132] = 1.0;
 sq1_lenEnable[133] = 1.0;
 sq1_lenEnable[134] = 1.0;
 sq1_lenEnable[135] = 1.0;
 sq1_lenEnable[136] = 1.0;
 sq1_lenEnable[137] = 1.0;
 sq1_lenEnable[138] = 1.0;
 sq1_lenEnable[139] = 1.0;
 sq1_lenEnable[140] = 1.0;
 sq1_lenEnable[141] = 1.0;
 sq1_lenEnable[142] = 1.0;
 sq1_lenEnable[143] = 1.0;
 sq1_lenEnable[144] = 1.0;
 sq1_lenEnable[145] = 1.0;
 sq1_lenEnable[146] = 1.0;
 sq1_lenEnable[147] = 1.0;
 sq1_lenEnable[148] = 1.0;
 sq1_lenEnable[149] = 1.0;
 sq1_lenEnable[150] = 1.0;
 sq1_lenEnable[151] = 1.0;
 sq1_lenEnable[152] = 1.0;
 sq1_lenEnable[153] = 1.0;
 sq1_lenEnable[154] = 1.0;
 sq1_lenEnable[155] = 1.0;
 sq1_lenEnable[156] = 1.0;
 sq1_lenEnable[157] = 1.0;
 sq1_lenEnable[158] = 1.0;
 sq1_lenEnable[159] = 1.0;
 sq1_lenEnable[160] = 1.0;
 sq1_lenEnable[161] = 1.0;
 sq1_lenEnable[162] = 1.0;
 sq1_lenEnable[163] = 1.0;
 sq1_lenEnable[164] = 1.0;
 sq1_lenEnable[165] = 1.0;
 sq1_lenEnable[166] = 1.0;
 sq1_lenEnable[167] = 1.0;
 sq1_lenEnable[168] = 1.0;
 sq1_lenEnable[169] = 1.0;
 sq1_lenEnable[170] = 1.0;
 sq1_lenEnable[171] = 1.0;
 sq1_lenEnable[172] = 1.0;
 sq1_lenEnable[173] = 1.0;
 sq1_lenEnable[174] = 1.0;
 sq1_lenEnable[175] = 1.0;
 sq1_lenEnable[176] = 1.0;
 sq1_lenEnable[177] = 1.0;
 sq1_lenEnable[178] = 1.0;
 sq1_lenEnable[179] = 1.0;
 sq1_lenEnable[180] = 1.0;
 sq1_lenEnable[181] = 1.0;
 sq1_lenEnable[182] = 1.0;
 sq1_lenEnable[183] = 1.0;
 sq1_lenEnable[184] = 1.0;
 sq1_lenEnable[185] = 1.0;
 sq1_lenEnable[186] = 1.0;
 sq1_lenEnable[187] = 1.0;
 sq1_lenEnable[188] = 1.0;
 sq1_lenEnable[189] = 1.0;
 sq1_lenEnable[190] = 1.0;
 sq1_lenEnable[191] = 1.0;
 sq1_lenEnable[192] = 1.0;
 sq1_lenEnable[193] = 1.0;
 sq1_lenEnable[194] = 1.0;
 sq1_lenEnable[195] = 1.0;
 sq1_lenEnable[196] = 1.0;
 sq1_lenEnable[197] = 1.0;
 sq1_lenEnable[198] = 1.0;
 sq1_lenEnable[199] = 1.0;
 sq1_lenEnable[200] = 1.0;
 sq1_lenEnable[201] = 1.0;
 sq1_lenEnable[202] = 1.0;
 sq1_lenEnable[203] = 1.0;
 sq1_lenEnable[204] = 1.0;
 sq1_lenEnable[205] = 1.0;
 sq1_lenEnable[206] = 1.0;
 sq1_lenEnable[207] = 1.0;
 sq1_lenEnable[208] = 1.0;
 sq1_lenEnable[209] = 1.0;
 sq1_lenEnable[210] = 1.0;
 sq1_lenEnable[211] = 1.0;
 sq1_lenEnable[212] = 1.0;
 sq1_lenEnable[213] = 1.0;
 sq1_lenEnable[214] = 1.0;
 sq1_lenEnable[215] = 1.0;
 sq1_lenEnable[216] = 1.0;
 sq1_lenEnable[217] = 1.0;
 sq1_lenEnable[218] = 1.0;
 sq1_lenEnable[219] = 1.0;
 sq1_lenEnable[220] = 1.0;
 sq1_lenEnable[221] = 1.0;
 sq1_lenEnable[222] = 1.0;
 sq1_lenEnable[223] = 1.0;
 sq1_lenEnable[224] = 1.0;
 sq1_lenEnable[225] = 1.0;
 sq1_lenEnable[226] = 1.0;
 sq1_lenEnable[227] = 1.0;
 sq1_lenEnable[228] = 1.0;
 sq1_lenEnable[229] = 1.0;
 sq1_lenEnable[230] = 1.0;
 sq1_lenEnable[231] = 1.0;
 sq1_lenEnable[232] = 1.0;
 sq1_lenEnable[233] = 1.0;
 sq1_lenEnable[234] = 1.0;
 sq1_lenEnable[235] = 1.0;
 sq1_lenEnable[236] = 1.0;
 sq1_lenEnable[237] = 1.0;
 sq1_lenEnable[238] = 1.0;
 sq1_lenEnable[239] = 1.0;
 sq1_lenEnable[240] = 1.0;
 sq1_lenEnable[241] = 1.0;
 sq1_lenEnable[242] = 1.0;
 sq1_lenEnable[243] = 1.0;
 sq1_lenEnable[244] = 1.0;
 sq1_lenEnable[245] = 1.0;
 sq1_lenEnable[246] = 1.0;
 sq1_lenEnable[247] = 1.0;
 sq1_lenEnable[248] = 1.0;
 sq1_lenEnable[249] = 1.0;
 sq1_lenEnable[250] = 1.0;
 sq1_lenEnable[251] = 1.0;
 sq1_lenEnable[252] = 1.0;
 sq1_lenEnable[253] = 1.0;
 sq1_lenEnable[254] = 1.0;
 sq1_lenEnable[255] = 1.0;
 sq1_lenEnable[256] = 1.0;
 sq1_lenEnable[257] = 1.0;
 sq1_lenEnable[258] = 1.0;
 sq1_lenEnable[259] = 1.0;
 sq1_lenEnable[260] = 1.0;
 sq1_lenEnable[261] = 1.0;
 sq1_lenEnable[262] = 1.0;
 sq1_lenEnable[263] = 1.0;
 sq1_lenEnable[264] = 1.0;
 sq1_lenEnable[265] = 1.0;
 sq1_lenEnable[266] = 1.0;
 sq1_lenEnable[267] = 1.0;
 sq1_lenEnable[268] = 1.0;
 sq1_lenEnable[269] = 1.0;
 sq1_lenEnable[270] = 1.0;
 sq1_lenEnable[271] = 1.0;
 sq1_lenEnable[272] = 1.0;
 sq1_lenEnable[273] = 1.0;
 sq1_lenEnable[274] = 1.0;
 sq1_lenEnable[275] = 1.0;
 sq1_lenEnable[276] = 1.0;
 sq1_lenEnable[277] = 1.0;
 sq1_lenEnable[278] = 1.0;
 sq1_lenEnable[279] = 1.0;
 sq1_lenEnable[280] = 1.0;
 sq1_lenEnable[281] = 1.0;
 sq1_lenEnable[282] = 1.0;
 sq1_lenEnable[283] = 1.0;
 sq1_lenEnable[284] = 1.0;
 sq1_lenEnable[285] = 1.0;
 sq1_lenEnable[286] = 1.0;
 sq1_lenEnable[287] = 1.0;
 sq1_lenEnable[288] = 1.0;
 sq1_lenEnable[289] = 1.0;
 sq1_lenEnable[290] = 1.0;
 sq1_lenEnable[291] = 1.0;
 sq1_lenEnable[292] = 1.0;
 sq1_lenEnable[293] = 1.0;
 sq1_lenEnable[294] = 1.0;
 sq1_lenEnable[295] = 1.0;
 sq1_lenEnable[296] = 1.0;
 sq1_lenEnable[297] = 1.0;
 sq1_lenEnable[298] = 1.0;
 sq1_lenEnable[299] = 1.0;
 sq1_lenEnable[300] = 1.0;
 sq1_lenEnable[301] = 1.0;
 sq1_lenEnable[302] = 1.0;
 sq1_lenEnable[303] = 1.0;
 sq1_lenEnable[304] = 1.0;
 sq1_lenEnable[305] = 1.0;
 sq1_lenEnable[306] = 1.0;
 sq1_lenEnable[307] = 1.0;
 sq1_lenEnable[308] = 1.0;
 sq1_lenEnable[309] = 1.0;
 sq1_lenEnable[310] = 1.0;
 sq1_lenEnable[311] = 1.0;
 sq1_lenEnable[312] = 1.0;
 sq1_lenEnable[313] = 1.0;
 sq1_lenEnable[314] = 1.0;
 sq1_lenEnable[315] = 1.0;
 sq1_lenEnable[316] = 1.0;
 sq1_lenEnable[317] = 1.0;
 sq1_lenEnable[318] = 1.0;
 sq1_lenEnable[319] = 1.0;
 sq1_lenEnable[320] = 1.0;
 sq1_lenEnable[321] = 1.0;
 sq1_lenEnable[322] = 1.0;
 sq1_lenEnable[323] = 1.0;
 sq1_lenEnable[324] = 1.0;
 sq1_lenEnable[325] = 1.0;
 sq1_lenEnable[326] = 1.0;
 sq1_lenEnable[327] = 1.0;
 sq1_lenEnable[328] = 1.0;
 sq1_lenEnable[329] = 1.0;
 sq1_lenEnable[330] = 1.0;
 sq1_lenEnable[331] = 1.0;
 sq1_lenEnable[332] = 1.0;
 sq1_lenEnable[333] = 1.0;
 sq1_lenEnable[334] = 1.0;
 sq1_lenEnable[335] = 1.0;
 sq1_lenEnable[336] = 1.0;
 sq1_lenEnable[337] = 1.0;
 sq1_lenEnable[338] = 1.0;
 sq1_lenEnable[339] = 1.0;
 sq1_lenEnable[340] = 1.0;
 sq1_lenEnable[341] = 1.0;
 sq1_lenEnable[342] = 1.0;
 sq1_lenEnable[343] = 1.0;
 sq1_lenEnable[344] = 1.0;
 sq1_lenEnable[345] = 1.0;
 sq1_lenEnable[346] = 1.0;
 sq1_lenEnable[347] = 1.0;
 sq1_lenEnable[348] = 1.0;
 sq1_lenEnable[349] = 1.0;
 sq1_lenEnable[350] = 1.0;
 sq1_lenEnable[351] = 1.0;
 sq1_lenEnable[352] = 1.0;
 sq1_lenEnable[353] = 1.0;
 sq1_lenEnable[354] = 1.0;
 sq1_lenEnable[355] = 1.0;
 sq1_lenEnable[356] = 1.0;
 sq1_lenEnable[357] = 1.0;
 sq1_lenEnable[358] = 1.0;
 sq1_lenEnable[359] = 1.0;
 sq1_lenEnable[360] = 1.0;
 sq1_lenEnable[361] = 1.0;
 sq1_lenEnable[362] = 1.0;
 sq1_lenEnable[363] = 1.0;
 sq1_lenEnable[364] = 1.0;
 sq1_lenEnable[365] = 1.0;
 sq1_lenEnable[366] = 1.0;
 sq1_lenEnable[367] = 1.0;
 sq1_lenEnable[368] = 1.0;
 sq1_lenEnable[369] = 1.0;
 sq1_lenEnable[370] = 1.0;
 sq1_lenEnable[371] = 1.0;
 sq1_lenEnable[372] = 1.0;
 sq1_lenEnable[373] = 1.0;
 sq1_lenEnable[374] = 1.0;
 sq1_lenEnable[375] = 1.0;
 sq1_lenEnable[376] = 1.0;
 sq1_lenEnable[377] = 1.0;
 sq1_lenEnable[378] = 1.0;
 sq2_duty[0] = 2.0;
 sq2_duty[1] = 2.0;
 sq2_duty[2] = 2.0;
 sq2_duty[3] = 2.0;
 sq2_duty[4] = 2.0;
 sq2_duty[5] = 2.0;
 sq2_duty[6] = 2.0;
 sq2_duty[7] = 2.0;
 sq2_duty[8] = 2.0;
 sq2_duty[9] = 2.0;
 sq2_duty[10] = 2.0;
 sq2_duty[11] = 2.0;
 sq2_duty[12] = 2.0;
 sq2_duty[13] = 2.0;
 sq2_duty[14] = 2.0;
 sq2_duty[15] = 2.0;
 sq2_duty[16] = 2.0;
 sq2_duty[17] = 2.0;
 sq2_duty[18] = 2.0;
 sq2_duty[19] = 2.0;
 sq2_duty[20] = 2.0;
 sq2_duty[21] = 2.0;
 sq2_duty[22] = 2.0;
 sq2_duty[23] = 2.0;
 sq2_duty[24] = 2.0;
 sq2_duty[25] = 2.0;
 sq2_duty[26] = 2.0;
 sq2_duty[27] = 2.0;
 sq2_duty[28] = 2.0;
 sq2_duty[29] = 2.0;
 sq2_duty[30] = 2.0;
 sq2_duty[31] = 2.0;
 sq2_duty[32] = 2.0;
 sq2_duty[33] = 2.0;
 sq2_duty[34] = 2.0;
 sq2_duty[35] = 2.0;
 sq2_duty[36] = 2.0;
 sq2_duty[37] = 2.0;
 sq2_duty[38] = 2.0;
 sq2_duty[39] = 2.0;
 sq2_duty[40] = 2.0;
 sq2_duty[41] = 2.0;
 sq2_duty[42] = 2.0;
 sq2_duty[43] = 2.0;
 sq2_duty[44] = 2.0;
 sq2_duty[45] = 2.0;
 sq2_duty[46] = 2.0;
 sq2_duty[47] = 2.0;
 sq2_duty[48] = 2.0;
 sq2_duty[49] = 2.0;
 sq2_duty[50] = 2.0;
 sq2_duty[51] = 2.0;
 sq2_duty[52] = 2.0;
 sq2_duty[53] = 2.0;
 sq2_duty[54] = 2.0;
 sq2_duty[55] = 2.0;
 sq2_duty[56] = 2.0;
 sq2_duty[57] = 2.0;
 sq2_duty[58] = 2.0;
 sq2_duty[59] = 2.0;
 sq2_duty[60] = 2.0;
 sq2_duty[61] = 2.0;
 sq2_duty[62] = 2.0;
 sq2_duty[63] = 2.0;
 sq2_duty[64] = 2.0;
 sq2_duty[65] = 2.0;
 sq2_duty[66] = 2.0;
 sq2_duty[67] = 2.0;
 sq2_duty[68] = 2.0;
 sq2_duty[69] = 2.0;
 sq2_duty[70] = 2.0;
 sq2_duty[71] = 2.0;
 sq2_duty[72] = 2.0;
 sq2_duty[73] = 2.0;
 sq2_duty[74] = 2.0;
 sq2_duty[75] = 2.0;
 sq2_duty[76] = 2.0;
 sq2_duty[77] = 2.0;
 sq2_duty[78] = 2.0;
 sq2_duty[79] = 2.0;
 sq2_duty[80] = 2.0;
 sq2_duty[81] = 2.0;
 sq2_duty[82] = 2.0;
 sq2_duty[83] = 2.0;
 sq2_duty[84] = 2.0;
 sq2_duty[85] = 2.0;
 sq2_duty[86] = 2.0;
 sq2_duty[87] = 2.0;
 sq2_duty[88] = 2.0;
 sq2_duty[89] = 2.0;
 sq2_duty[90] = 2.0;
 sq2_duty[91] = 2.0;
 sq2_duty[92] = 2.0;
 sq2_duty[93] = 2.0;
 sq2_duty[94] = 2.0;
 sq2_duty[95] = 2.0;
 sq2_duty[96] = 2.0;
 sq2_duty[97] = 2.0;
 sq2_duty[98] = 2.0;
 sq2_duty[99] = 2.0;
 sq2_duty[100] = 2.0;
 sq2_duty[101] = 2.0;
 sq2_duty[102] = 2.0;
 sq2_duty[103] = 2.0;
 sq2_duty[104] = 2.0;
 sq2_duty[105] = 2.0;
 sq2_duty[106] = 2.0;
 sq2_duty[107] = 2.0;
 sq2_duty[108] = 2.0;
 sq2_duty[109] = 2.0;
 sq2_duty[110] = 2.0;
 sq2_duty[111] = 2.0;
 sq2_duty[112] = 2.0;
 sq2_duty[113] = 2.0;
 sq2_duty[114] = 2.0;
 sq2_duty[115] = 2.0;
 sq2_duty[116] = 2.0;
 sq2_duty[117] = 2.0;
 sq2_duty[118] = 2.0;
 sq2_duty[119] = 2.0;
 sq2_duty[120] = 2.0;
 sq2_duty[121] = 2.0;
 sq2_duty[122] = 2.0;
 sq2_duty[123] = 2.0;
 sq2_duty[124] = 2.0;
 sq2_duty[125] = 2.0;
 sq2_duty[126] = 2.0;
 sq2_duty[127] = 2.0;
 sq2_duty[128] = 2.0;
 sq2_duty[129] = 2.0;
 sq2_duty[130] = 2.0;
 sq2_duty[131] = 2.0;
 sq2_duty[132] = 2.0;
 sq2_duty[133] = 2.0;
 sq2_duty[134] = 2.0;
 sq2_duty[135] = 2.0;
 sq2_duty[136] = 2.0;
 sq2_duty[137] = 2.0;
 sq2_duty[138] = 2.0;
 sq2_duty[139] = 2.0;
 sq2_duty[140] = 2.0;
 sq2_duty[141] = 2.0;
 sq2_duty[142] = 2.0;
 sq2_duty[143] = 2.0;
 sq2_duty[144] = 2.0;
 sq2_duty[145] = 2.0;
 sq2_duty[146] = 2.0;
 sq2_duty[147] = 2.0;
 sq2_duty[148] = 2.0;
 sq2_duty[149] = 2.0;
 sq2_duty[150] = 2.0;
 sq2_duty[151] = 2.0;
 sq2_duty[152] = 2.0;
 sq2_duty[153] = 2.0;
 sq2_duty[154] = 2.0;
 sq2_duty[155] = 2.0;
 sq2_duty[156] = 2.0;
 sq2_duty[157] = 2.0;
 sq2_duty[158] = 2.0;
 sq2_duty[159] = 2.0;
 sq2_duty[160] = 2.0;
 sq2_duty[161] = 2.0;
 sq2_duty[162] = 2.0;
 sq2_duty[163] = 2.0;
 sq2_duty[164] = 2.0;
 sq2_duty[165] = 2.0;
 sq2_duty[166] = 2.0;
 sq2_duty[167] = 2.0;
 sq2_duty[168] = 2.0;
 sq2_duty[169] = 2.0;
 sq2_duty[170] = 2.0;
 sq2_duty[171] = 2.0;
 sq2_duty[172] = 2.0;
 sq2_duty[173] = 2.0;
 sq2_duty[174] = 2.0;
 sq2_duty[175] = 2.0;
 sq2_duty[176] = 2.0;
 sq2_duty[177] = 2.0;
 sq2_duty[178] = 2.0;
 sq2_duty[179] = 2.0;
 sq2_duty[180] = 2.0;
 sq2_duty[181] = 2.0;
 sq2_duty[182] = 2.0;
 sq2_duty[183] = 2.0;
 sq2_duty[184] = 2.0;
 sq2_duty[185] = 2.0;
 sq2_duty[186] = 2.0;
 sq2_duty[187] = 2.0;
 sq2_duty[188] = 2.0;
 sq2_duty[189] = 2.0;
 sq2_duty[190] = 2.0;
 sq2_duty[191] = 2.0;
 sq2_duty[192] = 2.0;
 sq2_duty[193] = 2.0;
 sq2_duty[194] = 2.0;
 sq2_duty[195] = 2.0;
 sq2_duty[196] = 2.0;
 sq2_duty[197] = 2.0;
 sq2_duty[198] = 2.0;
 sq2_duty[199] = 2.0;
 sq2_duty[200] = 2.0;
 sq2_duty[201] = 2.0;
 sq2_duty[202] = 2.0;
 sq2_duty[203] = 2.0;
 sq2_duty[204] = 2.0;
 sq2_duty[205] = 2.0;
 sq2_duty[206] = 2.0;
 sq2_duty[207] = 2.0;
 sq2_duty[208] = 2.0;
 sq2_duty[209] = 2.0;
 sq2_duty[210] = 2.0;
 sq2_duty[211] = 2.0;
 sq2_duty[212] = 2.0;
 sq2_duty[213] = 2.0;
 sq2_duty[214] = 2.0;
 sq2_duty[215] = 2.0;
 sq2_duty[216] = 2.0;
 sq2_duty[217] = 2.0;
 sq2_duty[218] = 2.0;
 sq2_duty[219] = 2.0;
 sq2_duty[220] = 2.0;
 sq2_duty[221] = 2.0;
 sq2_duty[222] = 2.0;
 sq2_duty[223] = 2.0;
 sq2_duty[224] = 2.0;
 sq2_duty[225] = 2.0;
 sq2_duty[226] = 2.0;
 sq2_duty[227] = 2.0;
 sq2_duty[228] = 2.0;
 sq2_duty[229] = 2.0;
 sq2_duty[230] = 2.0;
 sq2_duty[231] = 2.0;
 sq2_duty[232] = 2.0;
 sq2_duty[233] = 2.0;
 sq2_duty[234] = 2.0;
 sq2_duty[235] = 2.0;
 sq2_duty[236] = 2.0;
 sq2_duty[237] = 2.0;
 sq2_duty[238] = 2.0;
 sq2_duty[239] = 2.0;
 sq2_duty[240] = 2.0;
 sq2_duty[241] = 2.0;
 sq2_duty[242] = 2.0;
 sq2_duty[243] = 2.0;
 sq2_duty[244] = 2.0;
 sq2_duty[245] = 2.0;
 sq2_duty[246] = 2.0;
 sq2_duty[247] = 2.0;
 sq2_duty[248] = 2.0;
 sq2_duty[249] = 2.0;
 sq2_duty[250] = 2.0;
 sq2_duty[251] = 2.0;
 sq2_duty[252] = 2.0;
 sq2_duty[253] = 2.0;
 sq2_duty[254] = 2.0;
 sq2_duty[255] = 2.0;
 sq2_duty[256] = 2.0;
 sq2_duty[257] = 2.0;
 sq2_duty[258] = 2.0;
 sq2_duty[259] = 2.0;
 sq2_duty[260] = 2.0;
 sq2_duty[261] = 2.0;
 sq2_duty[262] = 2.0;
 sq2_duty[263] = 2.0;
 sq2_duty[264] = 2.0;
 sq2_duty[265] = 2.0;
 sq2_duty[266] = 2.0;
 sq2_duty[267] = 2.0;
 sq2_duty[268] = 2.0;
 sq2_duty[269] = 2.0;
 sq2_duty[270] = 2.0;
 sq2_duty[271] = 2.0;
 sq2_duty[272] = 2.0;
 sq2_duty[273] = 2.0;
 sq2_duty[274] = 2.0;
 sq2_duty[275] = 2.0;
 sq2_duty[276] = 2.0;
 sq2_duty[277] = 2.0;
 sq2_duty[278] = 2.0;
 sq2_duty[279] = 2.0;
 sq2_duty[280] = 2.0;
 sq2_duty[281] = 2.0;
 sq2_duty[282] = 2.0;
 sq2_duty[283] = 2.0;
 sq2_duty[284] = 2.0;
 sq2_duty[285] = 2.0;
 sq2_duty[286] = 2.0;
 sq2_duty[287] = 2.0;
 sq2_duty[288] = 2.0;
 sq2_duty[289] = 2.0;
 sq2_duty[290] = 2.0;
 sq2_duty[291] = 2.0;
 sq2_duty[292] = 2.0;
 sq2_duty[293] = 2.0;
 sq2_duty[294] = 2.0;
 sq2_duty[295] = 2.0;
 sq2_duty[296] = 2.0;
 sq2_duty[297] = 2.0;
 sq2_duty[298] = 2.0;
 sq2_duty[299] = 2.0;
 sq2_duty[300] = 2.0;
 sq2_duty[301] = 2.0;
 sq2_duty[302] = 2.0;
 sq2_duty[303] = 2.0;
 sq2_duty[304] = 2.0;
 sq2_duty[305] = 2.0;
 sq2_duty[306] = 2.0;
 sq2_duty[307] = 2.0;
 sq2_duty[308] = 2.0;
 sq2_duty[309] = 2.0;
 sq2_duty[310] = 2.0;
 sq2_duty[311] = 2.0;
 sq2_duty[312] = 2.0;
 sq2_duty[313] = 2.0;
 sq2_duty[314] = 2.0;
 sq2_duty[315] = 2.0;
 sq2_duty[316] = 2.0;
 sq2_duty[317] = 2.0;
 sq2_duty[318] = 2.0;
 sq2_duty[319] = 2.0;
 sq2_duty[320] = 2.0;
 sq2_duty[321] = 2.0;
 sq2_duty[322] = 2.0;
 sq2_duty[323] = 2.0;
 sq2_duty[324] = 2.0;
 sq2_duty[325] = 2.0;
 sq2_duty[326] = 2.0;
 sq2_duty[327] = 2.0;
 sq2_duty[328] = 2.0;
 sq2_duty[329] = 2.0;
 sq2_duty[330] = 2.0;
 sq2_duty[331] = 2.0;
 sq2_duty[332] = 2.0;
 sq2_duty[333] = 2.0;
 sq2_duty[334] = 2.0;
 sq2_duty[335] = 2.0;
 sq2_duty[336] = 2.0;
 sq2_duty[337] = 2.0;
 sq2_duty[338] = 2.0;
 sq2_duty[339] = 2.0;
 sq2_duty[340] = 2.0;
 sq2_duty[341] = 2.0;
 sq2_duty[342] = 2.0;
 sq2_duty[343] = 2.0;
 sq2_duty[344] = 2.0;
 sq2_duty[345] = 2.0;
 sq2_duty[346] = 2.0;
 sq2_duty[347] = 2.0;
 sq2_duty[348] = 2.0;
 sq2_duty[349] = 2.0;
 sq2_duty[350] = 2.0;
 sq2_duty[351] = 2.0;
 sq2_duty[352] = 2.0;
 sq2_duty[353] = 2.0;
 sq2_duty[354] = 2.0;
 sq2_duty[355] = 2.0;
 sq2_duty[356] = 2.0;
 sq2_duty[357] = 2.0;
 sq2_duty[358] = 2.0;
 sq2_duty[359] = 2.0;
 sq2_duty[360] = 2.0;
 sq2_duty[361] = 2.0;
 sq2_duty[362] = 2.0;
 sq2_duty[363] = 2.0;
 sq2_duty[364] = 2.0;
 sq2_duty[365] = 2.0;
 sq2_duty[366] = 2.0;
 sq2_duty[367] = 2.0;
 sq2_duty[368] = 2.0;
 sq2_duty[369] = 2.0;
 sq2_duty[370] = 2.0;
 sq2_duty[371] = 2.0;
 sq2_duty[372] = 2.0;
 sq2_duty[373] = 2.0;
 sq2_duty[374] = 2.0;
 sq2_duty[375] = 2.0;
 sq2_duty[376] = 2.0;
 sq2_duty[377] = 2.0;
 sq2_duty[378] = 2.0;
 sq2_lenLoad[0] = 32.0;
 sq2_lenLoad[1] = 32.0;
 sq2_lenLoad[2] = 32.0;
 sq2_lenLoad[3] = 32.0;
 sq2_lenLoad[4] = 32.0;
 sq2_lenLoad[5] = 32.0;
 sq2_lenLoad[6] = 32.0;
 sq2_lenLoad[7] = 32.0;
 sq2_lenLoad[8] = 32.0;
 sq2_lenLoad[9] = 32.0;
 sq2_lenLoad[10] = 32.0;
 sq2_lenLoad[11] = 32.0;
 sq2_lenLoad[12] = 32.0;
 sq2_lenLoad[13] = 32.0;
 sq2_lenLoad[14] = 32.0;
 sq2_lenLoad[15] = 32.0;
 sq2_lenLoad[16] = 32.0;
 sq2_lenLoad[17] = 32.0;
 sq2_lenLoad[18] = 32.0;
 sq2_lenLoad[19] = 32.0;
 sq2_lenLoad[20] = 32.0;
 sq2_lenLoad[21] = 32.0;
 sq2_lenLoad[22] = 32.0;
 sq2_lenLoad[23] = 32.0;
 sq2_lenLoad[24] = 32.0;
 sq2_lenLoad[25] = 32.0;
 sq2_lenLoad[26] = 32.0;
 sq2_lenLoad[27] = 32.0;
 sq2_lenLoad[28] = 32.0;
 sq2_lenLoad[29] = 32.0;
 sq2_lenLoad[30] = 32.0;
 sq2_lenLoad[31] = 32.0;
 sq2_lenLoad[32] = 32.0;
 sq2_lenLoad[33] = 32.0;
 sq2_lenLoad[34] = 32.0;
 sq2_lenLoad[35] = 32.0;
 sq2_lenLoad[36] = 32.0;
 sq2_lenLoad[37] = 32.0;
 sq2_lenLoad[38] = 32.0;
 sq2_lenLoad[39] = 32.0;
 sq2_lenLoad[40] = 32.0;
 sq2_lenLoad[41] = 32.0;
 sq2_lenLoad[42] = 32.0;
 sq2_lenLoad[43] = 32.0;
 sq2_lenLoad[44] = 32.0;
 sq2_lenLoad[45] = 32.0;
 sq2_lenLoad[46] = 32.0;
 sq2_lenLoad[47] = 32.0;
 sq2_lenLoad[48] = 32.0;
 sq2_lenLoad[49] = 32.0;
 sq2_lenLoad[50] = 32.0;
 sq2_lenLoad[51] = 32.0;
 sq2_lenLoad[52] = 32.0;
 sq2_lenLoad[53] = 32.0;
 sq2_lenLoad[54] = 32.0;
 sq2_lenLoad[55] = 32.0;
 sq2_lenLoad[56] = 32.0;
 sq2_lenLoad[57] = 32.0;
 sq2_lenLoad[58] = 32.0;
 sq2_lenLoad[59] = 32.0;
 sq2_lenLoad[60] = 32.0;
 sq2_lenLoad[61] = 32.0;
 sq2_lenLoad[62] = 32.0;
 sq2_lenLoad[63] = 32.0;
 sq2_lenLoad[64] = 32.0;
 sq2_lenLoad[65] = 32.0;
 sq2_lenLoad[66] = 32.0;
 sq2_lenLoad[67] = 32.0;
 sq2_lenLoad[68] = 32.0;
 sq2_lenLoad[69] = 32.0;
 sq2_lenLoad[70] = 32.0;
 sq2_lenLoad[71] = 32.0;
 sq2_lenLoad[72] = 32.0;
 sq2_lenLoad[73] = 32.0;
 sq2_lenLoad[74] = 32.0;
 sq2_lenLoad[75] = 32.0;
 sq2_lenLoad[76] = 32.0;
 sq2_lenLoad[77] = 32.0;
 sq2_lenLoad[78] = 32.0;
 sq2_lenLoad[79] = 32.0;
 sq2_lenLoad[80] = 32.0;
 sq2_lenLoad[81] = 32.0;
 sq2_lenLoad[82] = 32.0;
 sq2_lenLoad[83] = 32.0;
 sq2_lenLoad[84] = 32.0;
 sq2_lenLoad[85] = 32.0;
 sq2_lenLoad[86] = 32.0;
 sq2_lenLoad[87] = 32.0;
 sq2_lenLoad[88] = 32.0;
 sq2_lenLoad[89] = 32.0;
 sq2_lenLoad[90] = 32.0;
 sq2_lenLoad[91] = 32.0;
 sq2_lenLoad[92] = 32.0;
 sq2_lenLoad[93] = 32.0;
 sq2_lenLoad[94] = 32.0;
 sq2_lenLoad[95] = 32.0;
 sq2_lenLoad[96] = 32.0;
 sq2_lenLoad[97] = 32.0;
 sq2_lenLoad[98] = 32.0;
 sq2_lenLoad[99] = 32.0;
 sq2_lenLoad[100] = 32.0;
 sq2_lenLoad[101] = 32.0;
 sq2_lenLoad[102] = 32.0;
 sq2_lenLoad[103] = 32.0;
 sq2_lenLoad[104] = 32.0;
 sq2_lenLoad[105] = 32.0;
 sq2_lenLoad[106] = 32.0;
 sq2_lenLoad[107] = 32.0;
 sq2_lenLoad[108] = 32.0;
 sq2_lenLoad[109] = 32.0;
 sq2_lenLoad[110] = 32.0;
 sq2_lenLoad[111] = 32.0;
 sq2_lenLoad[112] = 32.0;
 sq2_lenLoad[113] = 32.0;
 sq2_lenLoad[114] = 32.0;
 sq2_lenLoad[115] = 32.0;
 sq2_lenLoad[116] = 32.0;
 sq2_lenLoad[117] = 32.0;
 sq2_lenLoad[118] = 32.0;
 sq2_lenLoad[119] = 32.0;
 sq2_lenLoad[120] = 32.0;
 sq2_lenLoad[121] = 32.0;
 sq2_lenLoad[122] = 32.0;
 sq2_lenLoad[123] = 32.0;
 sq2_lenLoad[124] = 32.0;
 sq2_lenLoad[125] = 32.0;
 sq2_lenLoad[126] = 32.0;
 sq2_lenLoad[127] = 32.0;
 sq2_lenLoad[128] = 32.0;
 sq2_lenLoad[129] = 32.0;
 sq2_lenLoad[130] = 32.0;
 sq2_lenLoad[131] = 32.0;
 sq2_lenLoad[132] = 32.0;
 sq2_lenLoad[133] = 32.0;
 sq2_lenLoad[134] = 32.0;
 sq2_lenLoad[135] = 32.0;
 sq2_lenLoad[136] = 32.0;
 sq2_lenLoad[137] = 32.0;
 sq2_lenLoad[138] = 32.0;
 sq2_lenLoad[139] = 32.0;
 sq2_lenLoad[140] = 32.0;
 sq2_lenLoad[141] = 32.0;
 sq2_lenLoad[142] = 32.0;
 sq2_lenLoad[143] = 32.0;
 sq2_lenLoad[144] = 32.0;
 sq2_lenLoad[145] = 32.0;
 sq2_lenLoad[146] = 32.0;
 sq2_lenLoad[147] = 32.0;
 sq2_lenLoad[148] = 32.0;
 sq2_lenLoad[149] = 32.0;
 sq2_lenLoad[150] = 32.0;
 sq2_lenLoad[151] = 32.0;
 sq2_lenLoad[152] = 32.0;
 sq2_lenLoad[153] = 32.0;
 sq2_lenLoad[154] = 32.0;
 sq2_lenLoad[155] = 32.0;
 sq2_lenLoad[156] = 32.0;
 sq2_lenLoad[157] = 32.0;
 sq2_lenLoad[158] = 32.0;
 sq2_lenLoad[159] = 32.0;
 sq2_lenLoad[160] = 32.0;
 sq2_lenLoad[161] = 32.0;
 sq2_lenLoad[162] = 32.0;
 sq2_lenLoad[163] = 32.0;
 sq2_lenLoad[164] = 32.0;
 sq2_lenLoad[165] = 32.0;
 sq2_lenLoad[166] = 32.0;
 sq2_lenLoad[167] = 32.0;
 sq2_lenLoad[168] = 32.0;
 sq2_lenLoad[169] = 32.0;
 sq2_lenLoad[170] = 32.0;
 sq2_lenLoad[171] = 32.0;
 sq2_lenLoad[172] = 32.0;
 sq2_lenLoad[173] = 32.0;
 sq2_lenLoad[174] = 32.0;
 sq2_lenLoad[175] = 32.0;
 sq2_lenLoad[176] = 32.0;
 sq2_lenLoad[177] = 32.0;
 sq2_lenLoad[178] = 32.0;
 sq2_lenLoad[179] = 32.0;
 sq2_lenLoad[180] = 32.0;
 sq2_lenLoad[181] = 32.0;
 sq2_lenLoad[182] = 32.0;
 sq2_lenLoad[183] = 32.0;
 sq2_lenLoad[184] = 32.0;
 sq2_lenLoad[185] = 32.0;
 sq2_lenLoad[186] = 32.0;
 sq2_lenLoad[187] = 32.0;
 sq2_lenLoad[188] = 32.0;
 sq2_lenLoad[189] = 32.0;
 sq2_lenLoad[190] = 32.0;
 sq2_lenLoad[191] = 32.0;
 sq2_lenLoad[192] = 32.0;
 sq2_lenLoad[193] = 32.0;
 sq2_lenLoad[194] = 32.0;
 sq2_lenLoad[195] = 32.0;
 sq2_lenLoad[196] = 32.0;
 sq2_lenLoad[197] = 32.0;
 sq2_lenLoad[198] = 32.0;
 sq2_lenLoad[199] = 32.0;
 sq2_lenLoad[200] = 32.0;
 sq2_lenLoad[201] = 32.0;
 sq2_lenLoad[202] = 32.0;
 sq2_lenLoad[203] = 32.0;
 sq2_lenLoad[204] = 32.0;
 sq2_lenLoad[205] = 32.0;
 sq2_lenLoad[206] = 32.0;
 sq2_lenLoad[207] = 32.0;
 sq2_lenLoad[208] = 32.0;
 sq2_lenLoad[209] = 32.0;
 sq2_lenLoad[210] = 32.0;
 sq2_lenLoad[211] = 32.0;
 sq2_lenLoad[212] = 32.0;
 sq2_lenLoad[213] = 32.0;
 sq2_lenLoad[214] = 32.0;
 sq2_lenLoad[215] = 32.0;
 sq2_lenLoad[216] = 32.0;
 sq2_lenLoad[217] = 32.0;
 sq2_lenLoad[218] = 32.0;
 sq2_lenLoad[219] = 32.0;
 sq2_lenLoad[220] = 32.0;
 sq2_lenLoad[221] = 32.0;
 sq2_lenLoad[222] = 32.0;
 sq2_lenLoad[223] = 32.0;
 sq2_lenLoad[224] = 32.0;
 sq2_lenLoad[225] = 32.0;
 sq2_lenLoad[226] = 32.0;
 sq2_lenLoad[227] = 32.0;
 sq2_lenLoad[228] = 32.0;
 sq2_lenLoad[229] = 32.0;
 sq2_lenLoad[230] = 32.0;
 sq2_lenLoad[231] = 32.0;
 sq2_lenLoad[232] = 32.0;
 sq2_lenLoad[233] = 32.0;
 sq2_lenLoad[234] = 32.0;
 sq2_lenLoad[235] = 32.0;
 sq2_lenLoad[236] = 32.0;
 sq2_lenLoad[237] = 32.0;
 sq2_lenLoad[238] = 32.0;
 sq2_lenLoad[239] = 32.0;
 sq2_lenLoad[240] = 32.0;
 sq2_lenLoad[241] = 32.0;
 sq2_lenLoad[242] = 32.0;
 sq2_lenLoad[243] = 32.0;
 sq2_lenLoad[244] = 32.0;
 sq2_lenLoad[245] = 32.0;
 sq2_lenLoad[246] = 32.0;
 sq2_lenLoad[247] = 32.0;
 sq2_lenLoad[248] = 32.0;
 sq2_lenLoad[249] = 32.0;
 sq2_lenLoad[250] = 32.0;
 sq2_lenLoad[251] = 32.0;
 sq2_lenLoad[252] = 32.0;
 sq2_lenLoad[253] = 32.0;
 sq2_lenLoad[254] = 32.0;
 sq2_lenLoad[255] = 32.0;
 sq2_lenLoad[256] = 32.0;
 sq2_lenLoad[257] = 32.0;
 sq2_lenLoad[258] = 32.0;
 sq2_lenLoad[259] = 32.0;
 sq2_lenLoad[260] = 32.0;
 sq2_lenLoad[261] = 32.0;
 sq2_lenLoad[262] = 32.0;
 sq2_lenLoad[263] = 32.0;
 sq2_lenLoad[264] = 32.0;
 sq2_lenLoad[265] = 32.0;
 sq2_lenLoad[266] = 32.0;
 sq2_lenLoad[267] = 32.0;
 sq2_lenLoad[268] = 32.0;
 sq2_lenLoad[269] = 32.0;
 sq2_lenLoad[270] = 32.0;
 sq2_lenLoad[271] = 32.0;
 sq2_lenLoad[272] = 32.0;
 sq2_lenLoad[273] = 32.0;
 sq2_lenLoad[274] = 32.0;
 sq2_lenLoad[275] = 32.0;
 sq2_lenLoad[276] = 32.0;
 sq2_lenLoad[277] = 32.0;
 sq2_lenLoad[278] = 32.0;
 sq2_lenLoad[279] = 32.0;
 sq2_lenLoad[280] = 32.0;
 sq2_lenLoad[281] = 32.0;
 sq2_lenLoad[282] = 32.0;
 sq2_lenLoad[283] = 32.0;
 sq2_lenLoad[284] = 32.0;
 sq2_lenLoad[285] = 32.0;
 sq2_lenLoad[286] = 32.0;
 sq2_lenLoad[287] = 32.0;
 sq2_lenLoad[288] = 32.0;
 sq2_lenLoad[289] = 32.0;
 sq2_lenLoad[290] = 32.0;
 sq2_lenLoad[291] = 32.0;
 sq2_lenLoad[292] = 32.0;
 sq2_lenLoad[293] = 32.0;
 sq2_lenLoad[294] = 32.0;
 sq2_lenLoad[295] = 32.0;
 sq2_lenLoad[296] = 32.0;
 sq2_lenLoad[297] = 32.0;
 sq2_lenLoad[298] = 32.0;
 sq2_lenLoad[299] = 32.0;
 sq2_lenLoad[300] = 32.0;
 sq2_lenLoad[301] = 32.0;
 sq2_lenLoad[302] = 32.0;
 sq2_lenLoad[303] = 32.0;
 sq2_lenLoad[304] = 32.0;
 sq2_lenLoad[305] = 32.0;
 sq2_lenLoad[306] = 32.0;
 sq2_lenLoad[307] = 32.0;
 sq2_lenLoad[308] = 32.0;
 sq2_lenLoad[309] = 32.0;
 sq2_lenLoad[310] = 32.0;
 sq2_lenLoad[311] = 32.0;
 sq2_lenLoad[312] = 32.0;
 sq2_lenLoad[313] = 32.0;
 sq2_lenLoad[314] = 32.0;
 sq2_lenLoad[315] = 32.0;
 sq2_lenLoad[316] = 32.0;
 sq2_lenLoad[317] = 32.0;
 sq2_lenLoad[318] = 32.0;
 sq2_lenLoad[319] = 32.0;
 sq2_lenLoad[320] = 32.0;
 sq2_lenLoad[321] = 32.0;
 sq2_lenLoad[322] = 32.0;
 sq2_lenLoad[323] = 32.0;
 sq2_lenLoad[324] = 32.0;
 sq2_lenLoad[325] = 32.0;
 sq2_lenLoad[326] = 32.0;
 sq2_lenLoad[327] = 32.0;
 sq2_lenLoad[328] = 32.0;
 sq2_lenLoad[329] = 32.0;
 sq2_lenLoad[330] = 32.0;
 sq2_lenLoad[331] = 32.0;
 sq2_lenLoad[332] = 32.0;
 sq2_lenLoad[333] = 32.0;
 sq2_lenLoad[334] = 32.0;
 sq2_lenLoad[335] = 32.0;
 sq2_lenLoad[336] = 32.0;
 sq2_lenLoad[337] = 32.0;
 sq2_lenLoad[338] = 32.0;
 sq2_lenLoad[339] = 32.0;
 sq2_lenLoad[340] = 32.0;
 sq2_lenLoad[341] = 32.0;
 sq2_lenLoad[342] = 32.0;
 sq2_lenLoad[343] = 32.0;
 sq2_lenLoad[344] = 32.0;
 sq2_lenLoad[345] = 32.0;
 sq2_lenLoad[346] = 32.0;
 sq2_lenLoad[347] = 32.0;
 sq2_lenLoad[348] = 32.0;
 sq2_lenLoad[349] = 32.0;
 sq2_lenLoad[350] = 32.0;
 sq2_lenLoad[351] = 32.0;
 sq2_lenLoad[352] = 32.0;
 sq2_lenLoad[353] = 32.0;
 sq2_lenLoad[354] = 32.0;
 sq2_lenLoad[355] = 32.0;
 sq2_lenLoad[356] = 32.0;
 sq2_lenLoad[357] = 32.0;
 sq2_lenLoad[358] = 32.0;
 sq2_lenLoad[359] = 32.0;
 sq2_lenLoad[360] = 32.0;
 sq2_lenLoad[361] = 32.0;
 sq2_lenLoad[362] = 32.0;
 sq2_lenLoad[363] = 32.0;
 sq2_lenLoad[364] = 32.0;
 sq2_lenLoad[365] = 32.0;
 sq2_lenLoad[366] = 32.0;
 sq2_lenLoad[367] = 32.0;
 sq2_lenLoad[368] = 32.0;
 sq2_lenLoad[369] = 32.0;
 sq2_lenLoad[370] = 32.0;
 sq2_lenLoad[371] = 32.0;
 sq2_lenLoad[372] = 32.0;
 sq2_lenLoad[373] = 32.0;
 sq2_lenLoad[374] = 32.0;
 sq2_lenLoad[375] = 32.0;
 sq2_lenLoad[376] = 32.0;
 sq2_lenLoad[377] = 32.0;
 sq2_lenLoad[378] = 32.0;
 sq2_startVol[0] = 12.0;
 sq2_startVol[1] = 12.0;
 sq2_startVol[2] = 12.0;
 sq2_startVol[3] = 12.0;
 sq2_startVol[4] = 12.0;
 sq2_startVol[5] = 12.0;
 sq2_startVol[6] = 12.0;
 sq2_startVol[7] = 12.0;
 sq2_startVol[8] = 12.0;
 sq2_startVol[9] = 12.0;
 sq2_startVol[10] = 12.0;
 sq2_startVol[11] = 12.0;
 sq2_startVol[12] = 12.0;
 sq2_startVol[13] = 12.0;
 sq2_startVol[14] = 12.0;
 sq2_startVol[15] = 12.0;
 sq2_startVol[16] = 12.0;
 sq2_startVol[17] = 12.0;
 sq2_startVol[18] = 12.0;
 sq2_startVol[19] = 12.0;
 sq2_startVol[20] = 12.0;
 sq2_startVol[21] = 12.0;
 sq2_startVol[22] = 12.0;
 sq2_startVol[23] = 12.0;
 sq2_startVol[24] = 12.0;
 sq2_startVol[25] = 12.0;
 sq2_startVol[26] = 12.0;
 sq2_startVol[27] = 12.0;
 sq2_startVol[28] = 12.0;
 sq2_startVol[29] = 12.0;
 sq2_startVol[30] = 12.0;
 sq2_startVol[31] = 12.0;
 sq2_startVol[32] = 12.0;
 sq2_startVol[33] = 12.0;
 sq2_startVol[34] = 12.0;
 sq2_startVol[35] = 12.0;
 sq2_startVol[36] = 12.0;
 sq2_startVol[37] = 12.0;
 sq2_startVol[38] = 12.0;
 sq2_startVol[39] = 12.0;
 sq2_startVol[40] = 12.0;
 sq2_startVol[41] = 12.0;
 sq2_startVol[42] = 12.0;
 sq2_startVol[43] = 12.0;
 sq2_startVol[44] = 12.0;
 sq2_startVol[45] = 12.0;
 sq2_startVol[46] = 12.0;
 sq2_startVol[47] = 12.0;
 sq2_startVol[48] = 12.0;
 sq2_startVol[49] = 12.0;
 sq2_startVol[50] = 12.0;
 sq2_startVol[51] = 12.0;
 sq2_startVol[52] = 12.0;
 sq2_startVol[53] = 12.0;
 sq2_startVol[54] = 12.0;
 sq2_startVol[55] = 12.0;
 sq2_startVol[56] = 12.0;
 sq2_startVol[57] = 12.0;
 sq2_startVol[58] = 12.0;
 sq2_startVol[59] = 12.0;
 sq2_startVol[60] = 12.0;
 sq2_startVol[61] = 12.0;
 sq2_startVol[62] = 12.0;
 sq2_startVol[63] = 12.0;
 sq2_startVol[64] = 12.0;
 sq2_startVol[65] = 12.0;
 sq2_startVol[66] = 12.0;
 sq2_startVol[67] = 12.0;
 sq2_startVol[68] = 12.0;
 sq2_startVol[69] = 12.0;
 sq2_startVol[70] = 12.0;
 sq2_startVol[71] = 12.0;
 sq2_startVol[72] = 12.0;
 sq2_startVol[73] = 12.0;
 sq2_startVol[74] = 12.0;
 sq2_startVol[75] = 12.0;
 sq2_startVol[76] = 12.0;
 sq2_startVol[77] = 12.0;
 sq2_startVol[78] = 12.0;
 sq2_startVol[79] = 12.0;
 sq2_startVol[80] = 12.0;
 sq2_startVol[81] = 12.0;
 sq2_startVol[82] = 12.0;
 sq2_startVol[83] = 12.0;
 sq2_startVol[84] = 12.0;
 sq2_startVol[85] = 12.0;
 sq2_startVol[86] = 12.0;
 sq2_startVol[87] = 12.0;
 sq2_startVol[88] = 12.0;
 sq2_startVol[89] = 12.0;
 sq2_startVol[90] = 12.0;
 sq2_startVol[91] = 12.0;
 sq2_startVol[92] = 12.0;
 sq2_startVol[93] = 12.0;
 sq2_startVol[94] = 12.0;
 sq2_startVol[95] = 12.0;
 sq2_startVol[96] = 12.0;
 sq2_startVol[97] = 12.0;
 sq2_startVol[98] = 12.0;
 sq2_startVol[99] = 12.0;
 sq2_startVol[100] = 12.0;
 sq2_startVol[101] = 12.0;
 sq2_startVol[102] = 12.0;
 sq2_startVol[103] = 12.0;
 sq2_startVol[104] = 12.0;
 sq2_startVol[105] = 12.0;
 sq2_startVol[106] = 12.0;
 sq2_startVol[107] = 12.0;
 sq2_startVol[108] = 12.0;
 sq2_startVol[109] = 12.0;
 sq2_startVol[110] = 12.0;
 sq2_startVol[111] = 12.0;
 sq2_startVol[112] = 12.0;
 sq2_startVol[113] = 12.0;
 sq2_startVol[114] = 12.0;
 sq2_startVol[115] = 12.0;
 sq2_startVol[116] = 12.0;
 sq2_startVol[117] = 12.0;
 sq2_startVol[118] = 12.0;
 sq2_startVol[119] = 12.0;
 sq2_startVol[120] = 12.0;
 sq2_startVol[121] = 12.0;
 sq2_startVol[122] = 12.0;
 sq2_startVol[123] = 12.0;
 sq2_startVol[124] = 12.0;
 sq2_startVol[125] = 12.0;
 sq2_startVol[126] = 12.0;
 sq2_startVol[127] = 12.0;
 sq2_startVol[128] = 12.0;
 sq2_startVol[129] = 12.0;
 sq2_startVol[130] = 12.0;
 sq2_startVol[131] = 12.0;
 sq2_startVol[132] = 12.0;
 sq2_startVol[133] = 12.0;
 sq2_startVol[134] = 12.0;
 sq2_startVol[135] = 12.0;
 sq2_startVol[136] = 12.0;
 sq2_startVol[137] = 12.0;
 sq2_startVol[138] = 12.0;
 sq2_startVol[139] = 12.0;
 sq2_startVol[140] = 12.0;
 sq2_startVol[141] = 12.0;
 sq2_startVol[142] = 12.0;
 sq2_startVol[143] = 12.0;
 sq2_startVol[144] = 12.0;
 sq2_startVol[145] = 12.0;
 sq2_startVol[146] = 12.0;
 sq2_startVol[147] = 12.0;
 sq2_startVol[148] = 12.0;
 sq2_startVol[149] = 12.0;
 sq2_startVol[150] = 12.0;
 sq2_startVol[151] = 12.0;
 sq2_startVol[152] = 12.0;
 sq2_startVol[153] = 12.0;
 sq2_startVol[154] = 12.0;
 sq2_startVol[155] = 12.0;
 sq2_startVol[156] = 12.0;
 sq2_startVol[157] = 12.0;
 sq2_startVol[158] = 12.0;
 sq2_startVol[159] = 12.0;
 sq2_startVol[160] = 12.0;
 sq2_startVol[161] = 12.0;
 sq2_startVol[162] = 12.0;
 sq2_startVol[163] = 12.0;
 sq2_startVol[164] = 12.0;
 sq2_startVol[165] = 12.0;
 sq2_startVol[166] = 12.0;
 sq2_startVol[167] = 12.0;
 sq2_startVol[168] = 12.0;
 sq2_startVol[169] = 12.0;
 sq2_startVol[170] = 12.0;
 sq2_startVol[171] = 12.0;
 sq2_startVol[172] = 12.0;
 sq2_startVol[173] = 12.0;
 sq2_startVol[174] = 12.0;
 sq2_startVol[175] = 12.0;
 sq2_startVol[176] = 12.0;
 sq2_startVol[177] = 12.0;
 sq2_startVol[178] = 12.0;
 sq2_startVol[179] = 12.0;
 sq2_startVol[180] = 12.0;
 sq2_startVol[181] = 12.0;
 sq2_startVol[182] = 12.0;
 sq2_startVol[183] = 12.0;
 sq2_startVol[184] = 12.0;
 sq2_startVol[185] = 12.0;
 sq2_startVol[186] = 12.0;
 sq2_startVol[187] = 12.0;
 sq2_startVol[188] = 12.0;
 sq2_startVol[189] = 12.0;
 sq2_startVol[190] = 12.0;
 sq2_startVol[191] = 12.0;
 sq2_startVol[192] = 12.0;
 sq2_startVol[193] = 12.0;
 sq2_startVol[194] = 12.0;
 sq2_startVol[195] = 12.0;
 sq2_startVol[196] = 12.0;
 sq2_startVol[197] = 12.0;
 sq2_startVol[198] = 12.0;
 sq2_startVol[199] = 12.0;
 sq2_startVol[200] = 12.0;
 sq2_startVol[201] = 12.0;
 sq2_startVol[202] = 12.0;
 sq2_startVol[203] = 12.0;
 sq2_startVol[204] = 12.0;
 sq2_startVol[205] = 12.0;
 sq2_startVol[206] = 12.0;
 sq2_startVol[207] = 12.0;
 sq2_startVol[208] = 12.0;
 sq2_startVol[209] = 12.0;
 sq2_startVol[210] = 12.0;
 sq2_startVol[211] = 12.0;
 sq2_startVol[212] = 12.0;
 sq2_startVol[213] = 12.0;
 sq2_startVol[214] = 12.0;
 sq2_startVol[215] = 12.0;
 sq2_startVol[216] = 12.0;
 sq2_startVol[217] = 12.0;
 sq2_startVol[218] = 12.0;
 sq2_startVol[219] = 12.0;
 sq2_startVol[220] = 12.0;
 sq2_startVol[221] = 12.0;
 sq2_startVol[222] = 12.0;
 sq2_startVol[223] = 12.0;
 sq2_startVol[224] = 12.0;
 sq2_startVol[225] = 12.0;
 sq2_startVol[226] = 12.0;
 sq2_startVol[227] = 12.0;
 sq2_startVol[228] = 12.0;
 sq2_startVol[229] = 12.0;
 sq2_startVol[230] = 12.0;
 sq2_startVol[231] = 12.0;
 sq2_startVol[232] = 12.0;
 sq2_startVol[233] = 12.0;
 sq2_startVol[234] = 12.0;
 sq2_startVol[235] = 12.0;
 sq2_startVol[236] = 12.0;
 sq2_startVol[237] = 12.0;
 sq2_startVol[238] = 12.0;
 sq2_startVol[239] = 12.0;
 sq2_startVol[240] = 12.0;
 sq2_startVol[241] = 12.0;
 sq2_startVol[242] = 12.0;
 sq2_startVol[243] = 12.0;
 sq2_startVol[244] = 12.0;
 sq2_startVol[245] = 12.0;
 sq2_startVol[246] = 12.0;
 sq2_startVol[247] = 12.0;
 sq2_startVol[248] = 12.0;
 sq2_startVol[249] = 12.0;
 sq2_startVol[250] = 12.0;
 sq2_startVol[251] = 12.0;
 sq2_startVol[252] = 12.0;
 sq2_startVol[253] = 12.0;
 sq2_startVol[254] = 12.0;
 sq2_startVol[255] = 12.0;
 sq2_startVol[256] = 12.0;
 sq2_startVol[257] = 12.0;
 sq2_startVol[258] = 12.0;
 sq2_startVol[259] = 12.0;
 sq2_startVol[260] = 12.0;
 sq2_startVol[261] = 12.0;
 sq2_startVol[262] = 12.0;
 sq2_startVol[263] = 12.0;
 sq2_startVol[264] = 12.0;
 sq2_startVol[265] = 12.0;
 sq2_startVol[266] = 12.0;
 sq2_startVol[267] = 12.0;
 sq2_startVol[268] = 12.0;
 sq2_startVol[269] = 12.0;
 sq2_startVol[270] = 12.0;
 sq2_startVol[271] = 12.0;
 sq2_startVol[272] = 12.0;
 sq2_startVol[273] = 12.0;
 sq2_startVol[274] = 12.0;
 sq2_startVol[275] = 12.0;
 sq2_startVol[276] = 12.0;
 sq2_startVol[277] = 12.0;
 sq2_startVol[278] = 12.0;
 sq2_startVol[279] = 12.0;
 sq2_startVol[280] = 12.0;
 sq2_startVol[281] = 12.0;
 sq2_startVol[282] = 12.0;
 sq2_startVol[283] = 12.0;
 sq2_startVol[284] = 12.0;
 sq2_startVol[285] = 12.0;
 sq2_startVol[286] = 12.0;
 sq2_startVol[287] = 12.0;
 sq2_startVol[288] = 12.0;
 sq2_startVol[289] = 12.0;
 sq2_startVol[290] = 12.0;
 sq2_startVol[291] = 12.0;
 sq2_startVol[292] = 12.0;
 sq2_startVol[293] = 12.0;
 sq2_startVol[294] = 12.0;
 sq2_startVol[295] = 12.0;
 sq2_startVol[296] = 12.0;
 sq2_startVol[297] = 12.0;
 sq2_startVol[298] = 12.0;
 sq2_startVol[299] = 12.0;
 sq2_startVol[300] = 12.0;
 sq2_startVol[301] = 12.0;
 sq2_startVol[302] = 12.0;
 sq2_startVol[303] = 12.0;
 sq2_startVol[304] = 12.0;
 sq2_startVol[305] = 12.0;
 sq2_startVol[306] = 12.0;
 sq2_startVol[307] = 12.0;
 sq2_startVol[308] = 12.0;
 sq2_startVol[309] = 12.0;
 sq2_startVol[310] = 12.0;
 sq2_startVol[311] = 12.0;
 sq2_startVol[312] = 12.0;
 sq2_startVol[313] = 12.0;
 sq2_startVol[314] = 12.0;
 sq2_startVol[315] = 12.0;
 sq2_startVol[316] = 12.0;
 sq2_startVol[317] = 12.0;
 sq2_startVol[318] = 12.0;
 sq2_startVol[319] = 12.0;
 sq2_startVol[320] = 12.0;
 sq2_startVol[321] = 12.0;
 sq2_startVol[322] = 12.0;
 sq2_startVol[323] = 12.0;
 sq2_startVol[324] = 12.0;
 sq2_startVol[325] = 12.0;
 sq2_startVol[326] = 12.0;
 sq2_startVol[327] = 12.0;
 sq2_startVol[328] = 12.0;
 sq2_startVol[329] = 12.0;
 sq2_startVol[330] = 12.0;
 sq2_startVol[331] = 12.0;
 sq2_startVol[332] = 12.0;
 sq2_startVol[333] = 12.0;
 sq2_startVol[334] = 12.0;
 sq2_startVol[335] = 12.0;
 sq2_startVol[336] = 12.0;
 sq2_startVol[337] = 12.0;
 sq2_startVol[338] = 12.0;
 sq2_startVol[339] = 12.0;
 sq2_startVol[340] = 12.0;
 sq2_startVol[341] = 12.0;
 sq2_startVol[342] = 12.0;
 sq2_startVol[343] = 12.0;
 sq2_startVol[344] = 12.0;
 sq2_startVol[345] = 12.0;
 sq2_startVol[346] = 12.0;
 sq2_startVol[347] = 12.0;
 sq2_startVol[348] = 12.0;
 sq2_startVol[349] = 12.0;
 sq2_startVol[350] = 12.0;
 sq2_startVol[351] = 12.0;
 sq2_startVol[352] = 12.0;
 sq2_startVol[353] = 12.0;
 sq2_startVol[354] = 12.0;
 sq2_startVol[355] = 12.0;
 sq2_startVol[356] = 12.0;
 sq2_startVol[357] = 12.0;
 sq2_startVol[358] = 12.0;
 sq2_startVol[359] = 12.0;
 sq2_startVol[360] = 12.0;
 sq2_startVol[361] = 12.0;
 sq2_startVol[362] = 12.0;
 sq2_startVol[363] = 12.0;
 sq2_startVol[364] = 12.0;
 sq2_startVol[365] = 12.0;
 sq2_startVol[366] = 12.0;
 sq2_startVol[367] = 12.0;
 sq2_startVol[368] = 12.0;
 sq2_startVol[369] = 12.0;
 sq2_startVol[370] = 12.0;
 sq2_startVol[371] = 12.0;
 sq2_startVol[372] = 12.0;
 sq2_startVol[373] = 12.0;
 sq2_startVol[374] = 12.0;
 sq2_startVol[375] = 12.0;
 sq2_startVol[376] = 12.0;
 sq2_startVol[377] = 12.0;
 sq2_startVol[378] = 12.0;
 sq2_envAdd[0] = 0.0;
 sq2_envAdd[1] = 0.0;
 sq2_envAdd[2] = 0.0;
 sq2_envAdd[3] = 0.0;
 sq2_envAdd[4] = 0.0;
 sq2_envAdd[5] = 0.0;
 sq2_envAdd[6] = 0.0;
 sq2_envAdd[7] = 0.0;
 sq2_envAdd[8] = 0.0;
 sq2_envAdd[9] = 0.0;
 sq2_envAdd[10] = 0.0;
 sq2_envAdd[11] = 0.0;
 sq2_envAdd[12] = 0.0;
 sq2_envAdd[13] = 0.0;
 sq2_envAdd[14] = 0.0;
 sq2_envAdd[15] = 0.0;
 sq2_envAdd[16] = 0.0;
 sq2_envAdd[17] = 0.0;
 sq2_envAdd[18] = 0.0;
 sq2_envAdd[19] = 0.0;
 sq2_envAdd[20] = 0.0;
 sq2_envAdd[21] = 0.0;
 sq2_envAdd[22] = 0.0;
 sq2_envAdd[23] = 0.0;
 sq2_envAdd[24] = 0.0;
 sq2_envAdd[25] = 0.0;
 sq2_envAdd[26] = 0.0;
 sq2_envAdd[27] = 0.0;
 sq2_envAdd[28] = 0.0;
 sq2_envAdd[29] = 0.0;
 sq2_envAdd[30] = 0.0;
 sq2_envAdd[31] = 0.0;
 sq2_envAdd[32] = 0.0;
 sq2_envAdd[33] = 0.0;
 sq2_envAdd[34] = 0.0;
 sq2_envAdd[35] = 0.0;
 sq2_envAdd[36] = 0.0;
 sq2_envAdd[37] = 0.0;
 sq2_envAdd[38] = 0.0;
 sq2_envAdd[39] = 0.0;
 sq2_envAdd[40] = 0.0;
 sq2_envAdd[41] = 0.0;
 sq2_envAdd[42] = 0.0;
 sq2_envAdd[43] = 0.0;
 sq2_envAdd[44] = 0.0;
 sq2_envAdd[45] = 0.0;
 sq2_envAdd[46] = 0.0;
 sq2_envAdd[47] = 0.0;
 sq2_envAdd[48] = 0.0;
 sq2_envAdd[49] = 0.0;
 sq2_envAdd[50] = 0.0;
 sq2_envAdd[51] = 0.0;
 sq2_envAdd[52] = 0.0;
 sq2_envAdd[53] = 0.0;
 sq2_envAdd[54] = 0.0;
 sq2_envAdd[55] = 0.0;
 sq2_envAdd[56] = 0.0;
 sq2_envAdd[57] = 0.0;
 sq2_envAdd[58] = 0.0;
 sq2_envAdd[59] = 0.0;
 sq2_envAdd[60] = 0.0;
 sq2_envAdd[61] = 0.0;
 sq2_envAdd[62] = 0.0;
 sq2_envAdd[63] = 0.0;
 sq2_envAdd[64] = 0.0;
 sq2_envAdd[65] = 0.0;
 sq2_envAdd[66] = 0.0;
 sq2_envAdd[67] = 0.0;
 sq2_envAdd[68] = 0.0;
 sq2_envAdd[69] = 0.0;
 sq2_envAdd[70] = 0.0;
 sq2_envAdd[71] = 0.0;
 sq2_envAdd[72] = 0.0;
 sq2_envAdd[73] = 0.0;
 sq2_envAdd[74] = 0.0;
 sq2_envAdd[75] = 0.0;
 sq2_envAdd[76] = 0.0;
 sq2_envAdd[77] = 0.0;
 sq2_envAdd[78] = 0.0;
 sq2_envAdd[79] = 0.0;
 sq2_envAdd[80] = 0.0;
 sq2_envAdd[81] = 0.0;
 sq2_envAdd[82] = 0.0;
 sq2_envAdd[83] = 0.0;
 sq2_envAdd[84] = 0.0;
 sq2_envAdd[85] = 0.0;
 sq2_envAdd[86] = 0.0;
 sq2_envAdd[87] = 0.0;
 sq2_envAdd[88] = 0.0;
 sq2_envAdd[89] = 0.0;
 sq2_envAdd[90] = 0.0;
 sq2_envAdd[91] = 0.0;
 sq2_envAdd[92] = 0.0;
 sq2_envAdd[93] = 0.0;
 sq2_envAdd[94] = 0.0;
 sq2_envAdd[95] = 0.0;
 sq2_envAdd[96] = 0.0;
 sq2_envAdd[97] = 0.0;
 sq2_envAdd[98] = 0.0;
 sq2_envAdd[99] = 0.0;
 sq2_envAdd[100] = 0.0;
 sq2_envAdd[101] = 0.0;
 sq2_envAdd[102] = 0.0;
 sq2_envAdd[103] = 0.0;
 sq2_envAdd[104] = 0.0;
 sq2_envAdd[105] = 0.0;
 sq2_envAdd[106] = 0.0;
 sq2_envAdd[107] = 0.0;
 sq2_envAdd[108] = 0.0;
 sq2_envAdd[109] = 0.0;
 sq2_envAdd[110] = 0.0;
 sq2_envAdd[111] = 0.0;
 sq2_envAdd[112] = 0.0;
 sq2_envAdd[113] = 0.0;
 sq2_envAdd[114] = 0.0;
 sq2_envAdd[115] = 0.0;
 sq2_envAdd[116] = 0.0;
 sq2_envAdd[117] = 0.0;
 sq2_envAdd[118] = 0.0;
 sq2_envAdd[119] = 0.0;
 sq2_envAdd[120] = 0.0;
 sq2_envAdd[121] = 0.0;
 sq2_envAdd[122] = 0.0;
 sq2_envAdd[123] = 0.0;
 sq2_envAdd[124] = 0.0;
 sq2_envAdd[125] = 0.0;
 sq2_envAdd[126] = 0.0;
 sq2_envAdd[127] = 0.0;
 sq2_envAdd[128] = 0.0;
 sq2_envAdd[129] = 0.0;
 sq2_envAdd[130] = 0.0;
 sq2_envAdd[131] = 0.0;
 sq2_envAdd[132] = 0.0;
 sq2_envAdd[133] = 0.0;
 sq2_envAdd[134] = 0.0;
 sq2_envAdd[135] = 0.0;
 sq2_envAdd[136] = 0.0;
 sq2_envAdd[137] = 0.0;
 sq2_envAdd[138] = 0.0;
 sq2_envAdd[139] = 0.0;
 sq2_envAdd[140] = 0.0;
 sq2_envAdd[141] = 0.0;
 sq2_envAdd[142] = 0.0;
 sq2_envAdd[143] = 0.0;
 sq2_envAdd[144] = 0.0;
 sq2_envAdd[145] = 0.0;
 sq2_envAdd[146] = 0.0;
 sq2_envAdd[147] = 0.0;
 sq2_envAdd[148] = 0.0;
 sq2_envAdd[149] = 0.0;
 sq2_envAdd[150] = 0.0;
 sq2_envAdd[151] = 0.0;
 sq2_envAdd[152] = 0.0;
 sq2_envAdd[153] = 0.0;
 sq2_envAdd[154] = 0.0;
 sq2_envAdd[155] = 0.0;
 sq2_envAdd[156] = 0.0;
 sq2_envAdd[157] = 0.0;
 sq2_envAdd[158] = 0.0;
 sq2_envAdd[159] = 0.0;
 sq2_envAdd[160] = 0.0;
 sq2_envAdd[161] = 0.0;
 sq2_envAdd[162] = 0.0;
 sq2_envAdd[163] = 0.0;
 sq2_envAdd[164] = 0.0;
 sq2_envAdd[165] = 0.0;
 sq2_envAdd[166] = 0.0;
 sq2_envAdd[167] = 0.0;
 sq2_envAdd[168] = 0.0;
 sq2_envAdd[169] = 0.0;
 sq2_envAdd[170] = 0.0;
 sq2_envAdd[171] = 0.0;
 sq2_envAdd[172] = 0.0;
 sq2_envAdd[173] = 0.0;
 sq2_envAdd[174] = 0.0;
 sq2_envAdd[175] = 0.0;
 sq2_envAdd[176] = 0.0;
 sq2_envAdd[177] = 0.0;
 sq2_envAdd[178] = 0.0;
 sq2_envAdd[179] = 0.0;
 sq2_envAdd[180] = 0.0;
 sq2_envAdd[181] = 0.0;
 sq2_envAdd[182] = 0.0;
 sq2_envAdd[183] = 0.0;
 sq2_envAdd[184] = 0.0;
 sq2_envAdd[185] = 0.0;
 sq2_envAdd[186] = 0.0;
 sq2_envAdd[187] = 0.0;
 sq2_envAdd[188] = 0.0;
 sq2_envAdd[189] = 0.0;
 sq2_envAdd[190] = 0.0;
 sq2_envAdd[191] = 0.0;
 sq2_envAdd[192] = 0.0;
 sq2_envAdd[193] = 0.0;
 sq2_envAdd[194] = 0.0;
 sq2_envAdd[195] = 0.0;
 sq2_envAdd[196] = 0.0;
 sq2_envAdd[197] = 0.0;
 sq2_envAdd[198] = 0.0;
 sq2_envAdd[199] = 0.0;
 sq2_envAdd[200] = 0.0;
 sq2_envAdd[201] = 0.0;
 sq2_envAdd[202] = 0.0;
 sq2_envAdd[203] = 0.0;
 sq2_envAdd[204] = 0.0;
 sq2_envAdd[205] = 0.0;
 sq2_envAdd[206] = 0.0;
 sq2_envAdd[207] = 0.0;
 sq2_envAdd[208] = 0.0;
 sq2_envAdd[209] = 0.0;
 sq2_envAdd[210] = 0.0;
 sq2_envAdd[211] = 0.0;
 sq2_envAdd[212] = 0.0;
 sq2_envAdd[213] = 0.0;
 sq2_envAdd[214] = 0.0;
 sq2_envAdd[215] = 0.0;
 sq2_envAdd[216] = 0.0;
 sq2_envAdd[217] = 0.0;
 sq2_envAdd[218] = 0.0;
 sq2_envAdd[219] = 0.0;
 sq2_envAdd[220] = 0.0;
 sq2_envAdd[221] = 0.0;
 sq2_envAdd[222] = 0.0;
 sq2_envAdd[223] = 0.0;
 sq2_envAdd[224] = 0.0;
 sq2_envAdd[225] = 0.0;
 sq2_envAdd[226] = 0.0;
 sq2_envAdd[227] = 0.0;
 sq2_envAdd[228] = 0.0;
 sq2_envAdd[229] = 0.0;
 sq2_envAdd[230] = 0.0;
 sq2_envAdd[231] = 0.0;
 sq2_envAdd[232] = 0.0;
 sq2_envAdd[233] = 0.0;
 sq2_envAdd[234] = 0.0;
 sq2_envAdd[235] = 0.0;
 sq2_envAdd[236] = 0.0;
 sq2_envAdd[237] = 0.0;
 sq2_envAdd[238] = 0.0;
 sq2_envAdd[239] = 0.0;
 sq2_envAdd[240] = 0.0;
 sq2_envAdd[241] = 0.0;
 sq2_envAdd[242] = 0.0;
 sq2_envAdd[243] = 0.0;
 sq2_envAdd[244] = 0.0;
 sq2_envAdd[245] = 0.0;
 sq2_envAdd[246] = 0.0;
 sq2_envAdd[247] = 0.0;
 sq2_envAdd[248] = 0.0;
 sq2_envAdd[249] = 0.0;
 sq2_envAdd[250] = 0.0;
 sq2_envAdd[251] = 0.0;
 sq2_envAdd[252] = 0.0;
 sq2_envAdd[253] = 0.0;
 sq2_envAdd[254] = 0.0;
 sq2_envAdd[255] = 0.0;
 sq2_envAdd[256] = 0.0;
 sq2_envAdd[257] = 0.0;
 sq2_envAdd[258] = 0.0;
 sq2_envAdd[259] = 0.0;
 sq2_envAdd[260] = 0.0;
 sq2_envAdd[261] = 0.0;
 sq2_envAdd[262] = 0.0;
 sq2_envAdd[263] = 0.0;
 sq2_envAdd[264] = 0.0;
 sq2_envAdd[265] = 0.0;
 sq2_envAdd[266] = 0.0;
 sq2_envAdd[267] = 0.0;
 sq2_envAdd[268] = 0.0;
 sq2_envAdd[269] = 0.0;
 sq2_envAdd[270] = 0.0;
 sq2_envAdd[271] = 0.0;
 sq2_envAdd[272] = 0.0;
 sq2_envAdd[273] = 0.0;
 sq2_envAdd[274] = 0.0;
 sq2_envAdd[275] = 0.0;
 sq2_envAdd[276] = 0.0;
 sq2_envAdd[277] = 0.0;
 sq2_envAdd[278] = 0.0;
 sq2_envAdd[279] = 0.0;
 sq2_envAdd[280] = 0.0;
 sq2_envAdd[281] = 0.0;
 sq2_envAdd[282] = 0.0;
 sq2_envAdd[283] = 0.0;
 sq2_envAdd[284] = 0.0;
 sq2_envAdd[285] = 0.0;
 sq2_envAdd[286] = 0.0;
 sq2_envAdd[287] = 0.0;
 sq2_envAdd[288] = 0.0;
 sq2_envAdd[289] = 0.0;
 sq2_envAdd[290] = 0.0;
 sq2_envAdd[291] = 0.0;
 sq2_envAdd[292] = 0.0;
 sq2_envAdd[293] = 0.0;
 sq2_envAdd[294] = 0.0;
 sq2_envAdd[295] = 0.0;
 sq2_envAdd[296] = 0.0;
 sq2_envAdd[297] = 0.0;
 sq2_envAdd[298] = 0.0;
 sq2_envAdd[299] = 0.0;
 sq2_envAdd[300] = 0.0;
 sq2_envAdd[301] = 0.0;
 sq2_envAdd[302] = 0.0;
 sq2_envAdd[303] = 0.0;
 sq2_envAdd[304] = 0.0;
 sq2_envAdd[305] = 0.0;
 sq2_envAdd[306] = 0.0;
 sq2_envAdd[307] = 0.0;
 sq2_envAdd[308] = 0.0;
 sq2_envAdd[309] = 0.0;
 sq2_envAdd[310] = 0.0;
 sq2_envAdd[311] = 0.0;
 sq2_envAdd[312] = 0.0;
 sq2_envAdd[313] = 0.0;
 sq2_envAdd[314] = 0.0;
 sq2_envAdd[315] = 0.0;
 sq2_envAdd[316] = 0.0;
 sq2_envAdd[317] = 0.0;
 sq2_envAdd[318] = 0.0;
 sq2_envAdd[319] = 0.0;
 sq2_envAdd[320] = 0.0;
 sq2_envAdd[321] = 0.0;
 sq2_envAdd[322] = 0.0;
 sq2_envAdd[323] = 0.0;
 sq2_envAdd[324] = 0.0;
 sq2_envAdd[325] = 0.0;
 sq2_envAdd[326] = 0.0;
 sq2_envAdd[327] = 0.0;
 sq2_envAdd[328] = 0.0;
 sq2_envAdd[329] = 0.0;
 sq2_envAdd[330] = 0.0;
 sq2_envAdd[331] = 0.0;
 sq2_envAdd[332] = 0.0;
 sq2_envAdd[333] = 0.0;
 sq2_envAdd[334] = 0.0;
 sq2_envAdd[335] = 0.0;
 sq2_envAdd[336] = 0.0;
 sq2_envAdd[337] = 0.0;
 sq2_envAdd[338] = 0.0;
 sq2_envAdd[339] = 0.0;
 sq2_envAdd[340] = 0.0;
 sq2_envAdd[341] = 0.0;
 sq2_envAdd[342] = 0.0;
 sq2_envAdd[343] = 0.0;
 sq2_envAdd[344] = 0.0;
 sq2_envAdd[345] = 0.0;
 sq2_envAdd[346] = 0.0;
 sq2_envAdd[347] = 0.0;
 sq2_envAdd[348] = 0.0;
 sq2_envAdd[349] = 0.0;
 sq2_envAdd[350] = 0.0;
 sq2_envAdd[351] = 0.0;
 sq2_envAdd[352] = 0.0;
 sq2_envAdd[353] = 0.0;
 sq2_envAdd[354] = 0.0;
 sq2_envAdd[355] = 0.0;
 sq2_envAdd[356] = 0.0;
 sq2_envAdd[357] = 0.0;
 sq2_envAdd[358] = 0.0;
 sq2_envAdd[359] = 0.0;
 sq2_envAdd[360] = 0.0;
 sq2_envAdd[361] = 0.0;
 sq2_envAdd[362] = 0.0;
 sq2_envAdd[363] = 0.0;
 sq2_envAdd[364] = 0.0;
 sq2_envAdd[365] = 0.0;
 sq2_envAdd[366] = 0.0;
 sq2_envAdd[367] = 0.0;
 sq2_envAdd[368] = 0.0;
 sq2_envAdd[369] = 0.0;
 sq2_envAdd[370] = 0.0;
 sq2_envAdd[371] = 0.0;
 sq2_envAdd[372] = 0.0;
 sq2_envAdd[373] = 0.0;
 sq2_envAdd[374] = 0.0;
 sq2_envAdd[375] = 0.0;
 sq2_envAdd[376] = 0.0;
 sq2_envAdd[377] = 0.0;
 sq2_envAdd[378] = 0.0;
 sq2_period[0] = 4.0;
 sq2_period[1] = 4.0;
 sq2_period[2] = 4.0;
 sq2_period[3] = 4.0;
 sq2_period[4] = 4.0;
 sq2_period[5] = 4.0;
 sq2_period[6] = 4.0;
 sq2_period[7] = 4.0;
 sq2_period[8] = 4.0;
 sq2_period[9] = 4.0;
 sq2_period[10] = 4.0;
 sq2_period[11] = 4.0;
 sq2_period[12] = 4.0;
 sq2_period[13] = 4.0;
 sq2_period[14] = 4.0;
 sq2_period[15] = 4.0;
 sq2_period[16] = 4.0;
 sq2_period[17] = 4.0;
 sq2_period[18] = 4.0;
 sq2_period[19] = 4.0;
 sq2_period[20] = 4.0;
 sq2_period[21] = 4.0;
 sq2_period[22] = 4.0;
 sq2_period[23] = 4.0;
 sq2_period[24] = 4.0;
 sq2_period[25] = 4.0;
 sq2_period[26] = 4.0;
 sq2_period[27] = 4.0;
 sq2_period[28] = 4.0;
 sq2_period[29] = 4.0;
 sq2_period[30] = 4.0;
 sq2_period[31] = 4.0;
 sq2_period[32] = 4.0;
 sq2_period[33] = 4.0;
 sq2_period[34] = 4.0;
 sq2_period[35] = 4.0;
 sq2_period[36] = 4.0;
 sq2_period[37] = 4.0;
 sq2_period[38] = 4.0;
 sq2_period[39] = 4.0;
 sq2_period[40] = 4.0;
 sq2_period[41] = 4.0;
 sq2_period[42] = 4.0;
 sq2_period[43] = 4.0;
 sq2_period[44] = 4.0;
 sq2_period[45] = 4.0;
 sq2_period[46] = 4.0;
 sq2_period[47] = 4.0;
 sq2_period[48] = 4.0;
 sq2_period[49] = 4.0;
 sq2_period[50] = 4.0;
 sq2_period[51] = 4.0;
 sq2_period[52] = 4.0;
 sq2_period[53] = 4.0;
 sq2_period[54] = 4.0;
 sq2_period[55] = 4.0;
 sq2_period[56] = 4.0;
 sq2_period[57] = 4.0;
 sq2_period[58] = 4.0;
 sq2_period[59] = 4.0;
 sq2_period[60] = 4.0;
 sq2_period[61] = 4.0;
 sq2_period[62] = 4.0;
 sq2_period[63] = 4.0;
 sq2_period[64] = 4.0;
 sq2_period[65] = 4.0;
 sq2_period[66] = 4.0;
 sq2_period[67] = 4.0;
 sq2_period[68] = 4.0;
 sq2_period[69] = 4.0;
 sq2_period[70] = 4.0;
 sq2_period[71] = 4.0;
 sq2_period[72] = 4.0;
 sq2_period[73] = 4.0;
 sq2_period[74] = 4.0;
 sq2_period[75] = 4.0;
 sq2_period[76] = 4.0;
 sq2_period[77] = 4.0;
 sq2_period[78] = 4.0;
 sq2_period[79] = 4.0;
 sq2_period[80] = 4.0;
 sq2_period[81] = 4.0;
 sq2_period[82] = 4.0;
 sq2_period[83] = 4.0;
 sq2_period[84] = 4.0;
 sq2_period[85] = 4.0;
 sq2_period[86] = 4.0;
 sq2_period[87] = 4.0;
 sq2_period[88] = 4.0;
 sq2_period[89] = 4.0;
 sq2_period[90] = 4.0;
 sq2_period[91] = 4.0;
 sq2_period[92] = 4.0;
 sq2_period[93] = 4.0;
 sq2_period[94] = 4.0;
 sq2_period[95] = 4.0;
 sq2_period[96] = 4.0;
 sq2_period[97] = 4.0;
 sq2_period[98] = 4.0;
 sq2_period[99] = 4.0;
 sq2_period[100] = 4.0;
 sq2_period[101] = 4.0;
 sq2_period[102] = 4.0;
 sq2_period[103] = 4.0;
 sq2_period[104] = 4.0;
 sq2_period[105] = 4.0;
 sq2_period[106] = 4.0;
 sq2_period[107] = 4.0;
 sq2_period[108] = 4.0;
 sq2_period[109] = 4.0;
 sq2_period[110] = 4.0;
 sq2_period[111] = 4.0;
 sq2_period[112] = 4.0;
 sq2_period[113] = 4.0;
 sq2_period[114] = 4.0;
 sq2_period[115] = 4.0;
 sq2_period[116] = 4.0;
 sq2_period[117] = 4.0;
 sq2_period[118] = 4.0;
 sq2_period[119] = 4.0;
 sq2_period[120] = 4.0;
 sq2_period[121] = 4.0;
 sq2_period[122] = 4.0;
 sq2_period[123] = 4.0;
 sq2_period[124] = 4.0;
 sq2_period[125] = 4.0;
 sq2_period[126] = 4.0;
 sq2_period[127] = 4.0;
 sq2_period[128] = 4.0;
 sq2_period[129] = 4.0;
 sq2_period[130] = 4.0;
 sq2_period[131] = 4.0;
 sq2_period[132] = 4.0;
 sq2_period[133] = 4.0;
 sq2_period[134] = 4.0;
 sq2_period[135] = 4.0;
 sq2_period[136] = 4.0;
 sq2_period[137] = 4.0;
 sq2_period[138] = 4.0;
 sq2_period[139] = 4.0;
 sq2_period[140] = 4.0;
 sq2_period[141] = 4.0;
 sq2_period[142] = 4.0;
 sq2_period[143] = 4.0;
 sq2_period[144] = 4.0;
 sq2_period[145] = 4.0;
 sq2_period[146] = 4.0;
 sq2_period[147] = 4.0;
 sq2_period[148] = 4.0;
 sq2_period[149] = 4.0;
 sq2_period[150] = 4.0;
 sq2_period[151] = 4.0;
 sq2_period[152] = 4.0;
 sq2_period[153] = 4.0;
 sq2_period[154] = 4.0;
 sq2_period[155] = 4.0;
 sq2_period[156] = 4.0;
 sq2_period[157] = 4.0;
 sq2_period[158] = 4.0;
 sq2_period[159] = 4.0;
 sq2_period[160] = 4.0;
 sq2_period[161] = 4.0;
 sq2_period[162] = 4.0;
 sq2_period[163] = 4.0;
 sq2_period[164] = 4.0;
 sq2_period[165] = 4.0;
 sq2_period[166] = 4.0;
 sq2_period[167] = 4.0;
 sq2_period[168] = 4.0;
 sq2_period[169] = 4.0;
 sq2_period[170] = 4.0;
 sq2_period[171] = 4.0;
 sq2_period[172] = 4.0;
 sq2_period[173] = 4.0;
 sq2_period[174] = 4.0;
 sq2_period[175] = 4.0;
 sq2_period[176] = 4.0;
 sq2_period[177] = 4.0;
 sq2_period[178] = 4.0;
 sq2_period[179] = 4.0;
 sq2_period[180] = 4.0;
 sq2_period[181] = 4.0;
 sq2_period[182] = 4.0;
 sq2_period[183] = 4.0;
 sq2_period[184] = 4.0;
 sq2_period[185] = 4.0;
 sq2_period[186] = 4.0;
 sq2_period[187] = 4.0;
 sq2_period[188] = 4.0;
 sq2_period[189] = 4.0;
 sq2_period[190] = 4.0;
 sq2_period[191] = 4.0;
 sq2_period[192] = 4.0;
 sq2_period[193] = 4.0;
 sq2_period[194] = 4.0;
 sq2_period[195] = 4.0;
 sq2_period[196] = 4.0;
 sq2_period[197] = 4.0;
 sq2_period[198] = 4.0;
 sq2_period[199] = 4.0;
 sq2_period[200] = 4.0;
 sq2_period[201] = 4.0;
 sq2_period[202] = 4.0;
 sq2_period[203] = 4.0;
 sq2_period[204] = 4.0;
 sq2_period[205] = 4.0;
 sq2_period[206] = 4.0;
 sq2_period[207] = 4.0;
 sq2_period[208] = 4.0;
 sq2_period[209] = 4.0;
 sq2_period[210] = 4.0;
 sq2_period[211] = 4.0;
 sq2_period[212] = 4.0;
 sq2_period[213] = 4.0;
 sq2_period[214] = 4.0;
 sq2_period[215] = 4.0;
 sq2_period[216] = 4.0;
 sq2_period[217] = 4.0;
 sq2_period[218] = 4.0;
 sq2_period[219] = 4.0;
 sq2_period[220] = 4.0;
 sq2_period[221] = 4.0;
 sq2_period[222] = 4.0;
 sq2_period[223] = 4.0;
 sq2_period[224] = 4.0;
 sq2_period[225] = 4.0;
 sq2_period[226] = 4.0;
 sq2_period[227] = 4.0;
 sq2_period[228] = 4.0;
 sq2_period[229] = 4.0;
 sq2_period[230] = 4.0;
 sq2_period[231] = 4.0;
 sq2_period[232] = 4.0;
 sq2_period[233] = 4.0;
 sq2_period[234] = 4.0;
 sq2_period[235] = 4.0;
 sq2_period[236] = 4.0;
 sq2_period[237] = 4.0;
 sq2_period[238] = 4.0;
 sq2_period[239] = 4.0;
 sq2_period[240] = 4.0;
 sq2_period[241] = 4.0;
 sq2_period[242] = 4.0;
 sq2_period[243] = 4.0;
 sq2_period[244] = 4.0;
 sq2_period[245] = 4.0;
 sq2_period[246] = 4.0;
 sq2_period[247] = 4.0;
 sq2_period[248] = 4.0;
 sq2_period[249] = 4.0;
 sq2_period[250] = 4.0;
 sq2_period[251] = 4.0;
 sq2_period[252] = 4.0;
 sq2_period[253] = 4.0;
 sq2_period[254] = 4.0;
 sq2_period[255] = 4.0;
 sq2_period[256] = 4.0;
 sq2_period[257] = 4.0;
 sq2_period[258] = 4.0;
 sq2_period[259] = 4.0;
 sq2_period[260] = 4.0;
 sq2_period[261] = 4.0;
 sq2_period[262] = 4.0;
 sq2_period[263] = 4.0;
 sq2_period[264] = 4.0;
 sq2_period[265] = 4.0;
 sq2_period[266] = 4.0;
 sq2_period[267] = 4.0;
 sq2_period[268] = 4.0;
 sq2_period[269] = 4.0;
 sq2_period[270] = 4.0;
 sq2_period[271] = 4.0;
 sq2_period[272] = 4.0;
 sq2_period[273] = 4.0;
 sq2_period[274] = 4.0;
 sq2_period[275] = 4.0;
 sq2_period[276] = 4.0;
 sq2_period[277] = 4.0;
 sq2_period[278] = 4.0;
 sq2_period[279] = 4.0;
 sq2_period[280] = 4.0;
 sq2_period[281] = 4.0;
 sq2_period[282] = 4.0;
 sq2_period[283] = 4.0;
 sq2_period[284] = 4.0;
 sq2_period[285] = 4.0;
 sq2_period[286] = 4.0;
 sq2_period[287] = 4.0;
 sq2_period[288] = 4.0;
 sq2_period[289] = 4.0;
 sq2_period[290] = 4.0;
 sq2_period[291] = 4.0;
 sq2_period[292] = 4.0;
 sq2_period[293] = 4.0;
 sq2_period[294] = 4.0;
 sq2_period[295] = 4.0;
 sq2_period[296] = 4.0;
 sq2_period[297] = 4.0;
 sq2_period[298] = 4.0;
 sq2_period[299] = 4.0;
 sq2_period[300] = 4.0;
 sq2_period[301] = 4.0;
 sq2_period[302] = 4.0;
 sq2_period[303] = 4.0;
 sq2_period[304] = 4.0;
 sq2_period[305] = 4.0;
 sq2_period[306] = 4.0;
 sq2_period[307] = 4.0;
 sq2_period[308] = 4.0;
 sq2_period[309] = 4.0;
 sq2_period[310] = 4.0;
 sq2_period[311] = 4.0;
 sq2_period[312] = 4.0;
 sq2_period[313] = 4.0;
 sq2_period[314] = 4.0;
 sq2_period[315] = 4.0;
 sq2_period[316] = 4.0;
 sq2_period[317] = 4.0;
 sq2_period[318] = 4.0;
 sq2_period[319] = 4.0;
 sq2_period[320] = 4.0;
 sq2_period[321] = 4.0;
 sq2_period[322] = 4.0;
 sq2_period[323] = 4.0;
 sq2_period[324] = 4.0;
 sq2_period[325] = 4.0;
 sq2_period[326] = 4.0;
 sq2_period[327] = 4.0;
 sq2_period[328] = 4.0;
 sq2_period[329] = 4.0;
 sq2_period[330] = 4.0;
 sq2_period[331] = 4.0;
 sq2_period[332] = 4.0;
 sq2_period[333] = 4.0;
 sq2_period[334] = 4.0;
 sq2_period[335] = 4.0;
 sq2_period[336] = 4.0;
 sq2_period[337] = 4.0;
 sq2_period[338] = 4.0;
 sq2_period[339] = 4.0;
 sq2_period[340] = 4.0;
 sq2_period[341] = 4.0;
 sq2_period[342] = 4.0;
 sq2_period[343] = 4.0;
 sq2_period[344] = 4.0;
 sq2_period[345] = 4.0;
 sq2_period[346] = 4.0;
 sq2_period[347] = 4.0;
 sq2_period[348] = 4.0;
 sq2_period[349] = 4.0;
 sq2_period[350] = 4.0;
 sq2_period[351] = 4.0;
 sq2_period[352] = 4.0;
 sq2_period[353] = 4.0;
 sq2_period[354] = 4.0;
 sq2_period[355] = 4.0;
 sq2_period[356] = 4.0;
 sq2_period[357] = 4.0;
 sq2_period[358] = 4.0;
 sq2_period[359] = 4.0;
 sq2_period[360] = 4.0;
 sq2_period[361] = 4.0;
 sq2_period[362] = 4.0;
 sq2_period[363] = 4.0;
 sq2_period[364] = 4.0;
 sq2_period[365] = 4.0;
 sq2_period[366] = 4.0;
 sq2_period[367] = 4.0;
 sq2_period[368] = 4.0;
 sq2_period[369] = 4.0;
 sq2_period[370] = 4.0;
 sq2_period[371] = 4.0;
 sq2_period[372] = 4.0;
 sq2_period[373] = 4.0;
 sq2_period[374] = 4.0;
 sq2_period[375] = 4.0;
 sq2_period[376] = 4.0;
 sq2_period[377] = 4.0;
 sq2_period[378] = 4.0;
 sq2_freq[0] = 1517;
 sq2_freq[1] = 1517;
 sq2_freq[2] = 1517;
 sq2_freq[3] = 1517;
 sq2_freq[4] = 1517;
 sq2_freq[5] = 1517;
 sq2_freq[6] = 1517;
 sq2_freq[7] = 1517;
 sq2_freq[8] = 1517;
 sq2_freq[9] = 1517;
 sq2_freq[10] = 1517;
 sq2_freq[11] = 1517;
 sq2_freq[12] = 1517;
 sq2_freq[13] = 1517;
 sq2_freq[14] = 1517;
 sq2_freq[15] = 1517;
 sq2_freq[16] = 1517;
 sq2_freq[17] = 1517;
 sq2_freq[18] = 1517;
 sq2_freq[19] = 1517;
 sq2_freq[20] = 1452;
 sq2_freq[21] = 1452;
 sq2_freq[22] = 1452;
 sq2_freq[23] = 1452;
 sq2_freq[24] = 1517;
 sq2_freq[25] = 1517;
 sq2_freq[26] = 1517;
 sq2_freq[27] = 1517;
 sq2_freq[28] = 1517;
 sq2_freq[29] = 1517;
 sq2_freq[30] = 1517;
 sq2_freq[31] = 1517;
 sq2_freq[32] = 1517;
 sq2_freq[33] = 1517;
 sq2_freq[34] = 1517;
 sq2_freq[35] = 1517;
 sq2_freq[36] = 1517;
 sq2_freq[37] = 1517;
 sq2_freq[38] = 1517;
 sq2_freq[39] = 1546;
 sq2_freq[40] = 1546;
 sq2_freq[41] = 1546;
 sq2_freq[42] = 1602;
 sq2_freq[43] = 1602;
 sq2_freq[44] = 1602;
 sq2_freq[45] = 1650;
 sq2_freq[46] = 1650;
 sq2_freq[47] = 1650;
 sq2_freq[48] = 1673;
 sq2_freq[49] = 1673;
 sq2_freq[50] = 1673;
 sq2_freq[51] = 1673;
 sq2_freq[52] = 1673;
 sq2_freq[53] = 1673;
 sq2_freq[54] = 1714;
 sq2_freq[55] = 1714;
 sq2_freq[56] = 1714;
 sq2_freq[57] = 1714;
 sq2_freq[58] = 1714;
 sq2_freq[59] = 1714;
 sq2_freq[60] = 1714;
 sq2_freq[61] = 1714;
 sq2_freq[62] = 1714;
 sq2_freq[63] = 1750;
 sq2_freq[64] = 1750;
 sq2_freq[65] = 1750;
 sq2_freq[66] = 1783;
 sq2_freq[67] = 1783;
 sq2_freq[68] = 1783;
 sq2_freq[69] = 1798;
 sq2_freq[70] = 1798;
 sq2_freq[71] = 1798;
 sq2_freq[72] = 1825;
 sq2_freq[73] = 1825;
 sq2_freq[74] = 1825;
 sq2_freq[75] = 1825;
 sq2_freq[76] = 1825;
 sq2_freq[77] = 1825;
 sq2_freq[78] = 1825;
 sq2_freq[79] = 1825;
 sq2_freq[80] = 1825;
 sq2_freq[81] = 1825;
 sq2_freq[82] = 1825;
 sq2_freq[83] = 1825;
 sq2_freq[84] = 1673;
 sq2_freq[85] = 1673;
 sq2_freq[86] = 1673;
 sq2_freq[87] = 1673;
 sq2_freq[88] = 1714;
 sq2_freq[89] = 1714;
 sq2_freq[90] = 1714;
 sq2_freq[91] = 1714;
 sq2_freq[92] = 1750;
 sq2_freq[93] = 1750;
 sq2_freq[94] = 1750;
 sq2_freq[95] = 1750;
 sq2_freq[96] = 1627;
 sq2_freq[97] = 1627;
 sq2_freq[98] = 1627;
 sq2_freq[99] = 1627;
 sq2_freq[100] = 1627;
 sq2_freq[101] = 1627;
 sq2_freq[102] = 1627;
 sq2_freq[103] = 1627;
 sq2_freq[104] = 1627;
 sq2_freq[105] = 1627;
 sq2_freq[106] = 1627;
 sq2_freq[107] = 1627;
 sq2_freq[108] = 1627;
 sq2_freq[109] = 1627;
 sq2_freq[110] = 1627;
 sq2_freq[111] = 1673;
 sq2_freq[112] = 1673;
 sq2_freq[113] = 1673;
 sq2_freq[114] = 1714;
 sq2_freq[115] = 1714;
 sq2_freq[116] = 1714;
 sq2_freq[117] = 1750;
 sq2_freq[118] = 1750;
 sq2_freq[119] = 1750;
 sq2_freq[120] = 1767;
 sq2_freq[121] = 1767;
 sq2_freq[122] = 1767;
 sq2_freq[123] = 1767;
 sq2_freq[124] = 1767;
 sq2_freq[125] = 1767;
 sq2_freq[126] = 1767;
 sq2_freq[127] = 1767;
 sq2_freq[128] = 1767;
 sq2_freq[129] = 1767;
 sq2_freq[130] = 1767;
 sq2_freq[131] = 1767;
 sq2_freq[132] = 1767;
 sq2_freq[133] = 1767;
 sq2_freq[134] = 1767;
 sq2_freq[135] = 1767;
 sq2_freq[136] = 1750;
 sq2_freq[137] = 1750;
 sq2_freq[138] = 1750;
 sq2_freq[139] = 1750;
 sq2_freq[140] = 1714;
 sq2_freq[141] = 1714;
 sq2_freq[142] = 1714;
 sq2_freq[143] = 1714;
 sq2_freq[144] = 1767;
 sq2_freq[145] = 1767;
 sq2_freq[146] = 1767;
 sq2_freq[147] = 1767;
 sq2_freq[148] = 1767;
 sq2_freq[149] = 1767;
 sq2_freq[150] = 1767;
 sq2_freq[151] = 1767;
 sq2_freq[152] = 1714;
 sq2_freq[153] = 1714;
 sq2_freq[154] = 1714;
 sq2_freq[155] = 1714;
 sq2_freq[156] = 1673;
 sq2_freq[157] = 1673;
 sq2_freq[158] = 1673;
 sq2_freq[159] = 1673;
 sq2_freq[160] = 1673;
 sq2_freq[161] = 1673;
 sq2_freq[162] = 1673;
 sq2_freq[163] = 1673;
 sq2_freq[164] = 1627;
 sq2_freq[165] = 1627;
 sq2_freq[166] = 1627;
 sq2_freq[167] = 1627;
 sq2_freq[168] = 1673;
 sq2_freq[169] = 1673;
 sq2_freq[170] = 1673;
 sq2_freq[171] = 1673;
 sq2_freq[172] = 1673;
 sq2_freq[173] = 1673;
 sq2_freq[174] = 1673;
 sq2_freq[175] = 1673;
 sq2_freq[176] = 1673;
 sq2_freq[177] = 1673;
 sq2_freq[178] = 1673;
 sq2_freq[179] = 1673;
 sq2_freq[180] = 1673;
 sq2_freq[181] = 1673;
 sq2_freq[182] = 1673;
 sq2_freq[183] = 1673;
 sq2_freq[184] = 1627;
 sq2_freq[185] = 1627;
 sq2_freq[186] = 1627;
 sq2_freq[187] = 1627;
 sq2_freq[188] = 1673;
 sq2_freq[189] = 1673;
 sq2_freq[190] = 1673;
 sq2_freq[191] = 1673;
 sq2_freq[192] = 1627;
 sq2_freq[193] = 1627;
 sq2_freq[194] = 1627;
 sq2_freq[195] = 1627;
 sq2_freq[196] = 1627;
 sq2_freq[197] = 1627;
 sq2_freq[198] = 1627;
 sq2_freq[199] = 1627;
 sq2_freq[200] = 1627;
 sq2_freq[201] = 1602;
 sq2_freq[202] = 1602;
 sq2_freq[203] = 1602;
 sq2_freq[204] = 1627;
 sq2_freq[205] = 1627;
 sq2_freq[206] = 1627;
 sq2_freq[207] = 1627;
 sq2_freq[208] = 1627;
 sq2_freq[209] = 1627;
 sq2_freq[210] = 1627;
 sq2_freq[211] = 1627;
 sq2_freq[212] = 1627;
 sq2_freq[213] = 1673;
 sq2_freq[214] = 1673;
 sq2_freq[215] = 1673;
 sq2_freq[216] = 1714;
 sq2_freq[217] = 1714;
 sq2_freq[218] = 1714;
 sq2_freq[219] = 1714;
 sq2_freq[220] = 1714;
 sq2_freq[221] = 1714;
 sq2_freq[222] = 1714;
 sq2_freq[223] = 1714;
 sq2_freq[224] = 1714;
 sq2_freq[225] = 1714;
 sq2_freq[226] = 1714;
 sq2_freq[227] = 1714;
 sq2_freq[228] = 1673;
 sq2_freq[229] = 1673;
 sq2_freq[230] = 1673;
 sq2_freq[231] = 1673;
 sq2_freq[232] = 1673;
 sq2_freq[233] = 1673;
 sq2_freq[234] = 1627;
 sq2_freq[235] = 1627;
 sq2_freq[236] = 1627;
 sq2_freq[237] = 1627;
 sq2_freq[238] = 1627;
 sq2_freq[239] = 1627;
 sq2_freq[240] = 1602;
 sq2_freq[241] = 1602;
 sq2_freq[242] = 1602;
 sq2_freq[243] = 1602;
 sq2_freq[244] = 1602;
 sq2_freq[245] = 1602;
 sq2_freq[246] = 1602;
 sq2_freq[247] = 1602;
 sq2_freq[248] = 1602;
 sq2_freq[249] = 1546;
 sq2_freq[250] = 1546;
 sq2_freq[251] = 1546;
 sq2_freq[252] = 1602;
 sq2_freq[253] = 1602;
 sq2_freq[254] = 1602;
 sq2_freq[255] = 1602;
 sq2_freq[256] = 1602;
 sq2_freq[257] = 1602;
 sq2_freq[258] = 1602;
 sq2_freq[259] = 1602;
 sq2_freq[260] = 1602;
 sq2_freq[261] = 1627;
 sq2_freq[262] = 1627;
 sq2_freq[263] = 1627;
 sq2_freq[264] = 1673;
 sq2_freq[265] = 1673;
 sq2_freq[266] = 1673;
 sq2_freq[267] = 1673;
 sq2_freq[268] = 1673;
 sq2_freq[269] = 1673;
 sq2_freq[270] = 1673;
 sq2_freq[271] = 1673;
 sq2_freq[272] = 1673;
 sq2_freq[273] = 1673;
 sq2_freq[274] = 1673;
 sq2_freq[275] = 1673;
 sq2_freq[276] = 1627;
 sq2_freq[277] = 1627;
 sq2_freq[278] = 1627;
 sq2_freq[279] = 1627;
 sq2_freq[280] = 1627;
 sq2_freq[281] = 1627;
 sq2_freq[282] = 1602;
 sq2_freq[283] = 1602;
 sq2_freq[284] = 1602;
 sq2_freq[285] = 1602;
 sq2_freq[286] = 1602;
 sq2_freq[287] = 1602;
 sq2_freq[288] = 1575;
 sq2_freq[289] = 1575;
 sq2_freq[290] = 1575;
 sq2_freq[291] = 1575;
 sq2_freq[292] = 1575;
 sq2_freq[293] = 1575;
 sq2_freq[294] = 1575;
 sq2_freq[295] = 1575;
 sq2_freq[296] = 1575;
 sq2_freq[297] = 1575;
 sq2_freq[298] = 1575;
 sq2_freq[299] = 1575;
 sq2_freq[300] = 1575;
 sq2_freq[301] = 1575;
 sq2_freq[302] = 1575;
 sq2_freq[303] = 1575;
 sq2_freq[304] = 1575;
 sq2_freq[305] = 1575;
 sq2_freq[306] = 1575;
 sq2_freq[307] = 1575;
 sq2_freq[308] = 1575;
 sq2_freq[309] = 1602;
 sq2_freq[310] = 1602;
 sq2_freq[311] = 1602;
 sq2_freq[312] = 1650;
 sq2_freq[313] = 1650;
 sq2_freq[314] = 1650;
 sq2_freq[315] = 1650;
 sq2_freq[316] = 1650;
 sq2_freq[317] = 1650;
 sq2_freq[318] = 1650;
 sq2_freq[319] = 1650;
 sq2_freq[320] = 1650;
 sq2_freq[321] = 1694;
 sq2_freq[322] = 1694;
 sq2_freq[323] = 1694;
 sq2_freq[324] = 1714;
 sq2_freq[325] = 1714;
 sq2_freq[326] = 1714;
 sq2_freq[327] = 1714;
 sq2_freq[328] = 1714;
 sq2_freq[329] = 1714;
 sq2_freq[330] = 1750;
 sq2_freq[331] = 1750;
 sq2_freq[332] = 1750;
 sq2_freq[333] = 1750;
 sq2_freq[334] = 1750;
 sq2_freq[335] = 1750;
 sq2_freq[336] = 1602;
 sq2_freq[337] = 1602;
 sq2_freq[338] = 1602;
 sq2_freq[339] = 1602;
 sq2_freq[340] = 1602;
 sq2_freq[341] = 1602;
 sq2_freq[342] = 1602;
 sq2_freq[343] = 1602;
 sq2_freq[344] = 1602;
 sq2_freq[345] = 1602;
 sq2_freq[346] = 1602;
 sq2_freq[347] = 1602;
 sq2_freq[348] = 1602;
 sq2_freq[349] = 1602;
 sq2_freq[350] = 1602;
 sq2_freq[351] = 1602;
 sq2_freq[352] = 1602;
 sq2_freq[353] = 1602;
 sq2_freq[354] = 1602;
 sq2_freq[355] = 1602;
 sq2_freq[356] = 1602;
 sq2_freq[357] = 1602;
 sq2_freq[358] = 1602;
 sq2_freq[359] = 1602;
 sq2_freq[360] = 1602;
 sq2_freq[361] = 1602;
 sq2_freq[362] = 1602;
 sq2_freq[363] = 1602;
 sq2_freq[364] = 1602;
 sq2_freq[365] = 1602;
 sq2_freq[366] = 1602;
 sq2_freq[367] = 1602;
 sq2_freq[368] = 1602;
 sq2_freq[369] = 1602;
 sq2_freq[370] = 1602;
 sq2_freq[371] = 1602;
 sq2_freq[372] = 1602;
 sq2_freq[373] = 1602;
 sq2_freq[374] = 1602;
 sq2_freq[375] = 1602;
 sq2_freq[376] = 1602;
 sq2_freq[377] = 1602;
 sq2_freq[378] = 1602;
 sq2_trigger[0] = 1.0;
 sq2_trigger[1] = 0;
 sq2_trigger[2] = 0;
 sq2_trigger[3] = 0;
 sq2_trigger[4] = 0;
 sq2_trigger[5] = 0;
 sq2_trigger[6] = 0;
 sq2_trigger[7] = 0;
 sq2_trigger[8] = 0;
 sq2_trigger[9] = 0;
 sq2_trigger[10] = 0;
 sq2_trigger[11] = 0;
 sq2_trigger[12] = 1.0;
 sq2_trigger[13] = 0;
 sq2_trigger[14] = 0;
 sq2_trigger[15] = 0;
 sq2_trigger[16] = 1.0;
 sq2_trigger[17] = 0;
 sq2_trigger[18] = 0;
 sq2_trigger[19] = 0;
 sq2_trigger[20] = 1.0;
 sq2_trigger[21] = 0;
 sq2_trigger[22] = 0;
 sq2_trigger[23] = 0;
 sq2_trigger[24] = 1.0;
 sq2_trigger[25] = 0;
 sq2_trigger[26] = 0;
 sq2_trigger[27] = 0;
 sq2_trigger[28] = 0;
 sq2_trigger[29] = 0;
 sq2_trigger[30] = 0;
 sq2_trigger[31] = 0;
 sq2_trigger[32] = 0;
 sq2_trigger[33] = 0;
 sq2_trigger[34] = 0;
 sq2_trigger[35] = 0;
 sq2_trigger[36] = 1.0;
 sq2_trigger[37] = 0;
 sq2_trigger[38] = 0;
 sq2_trigger[39] = 1.0;
 sq2_trigger[40] = 0;
 sq2_trigger[41] = 0;
 sq2_trigger[42] = 1.0;
 sq2_trigger[43] = 0;
 sq2_trigger[44] = 0;
 sq2_trigger[45] = 1.0;
 sq2_trigger[46] = 0;
 sq2_trigger[47] = 0;
 sq2_trigger[48] = 1.0;
 sq2_trigger[49] = 0;
 sq2_trigger[50] = 0;
 sq2_trigger[51] = 0;
 sq2_trigger[52] = 0;
 sq2_trigger[53] = 0;
 sq2_trigger[54] = 1.0;
 sq2_trigger[55] = 0;
 sq2_trigger[56] = 0;
 sq2_trigger[57] = 0;
 sq2_trigger[58] = 0;
 sq2_trigger[59] = 0;
 sq2_trigger[60] = 1.0;
 sq2_trigger[61] = 0;
 sq2_trigger[62] = 0;
 sq2_trigger[63] = 1.0;
 sq2_trigger[64] = 0;
 sq2_trigger[65] = 0;
 sq2_trigger[66] = 1.0;
 sq2_trigger[67] = 0;
 sq2_trigger[68] = 0;
 sq2_trigger[69] = 1.0;
 sq2_trigger[70] = 0;
 sq2_trigger[71] = 0;
 sq2_trigger[72] = 1.0;
 sq2_trigger[73] = 0;
 sq2_trigger[74] = 0;
 sq2_trigger[75] = 0;
 sq2_trigger[76] = 0;
 sq2_trigger[77] = 0;
 sq2_trigger[78] = 0;
 sq2_trigger[79] = 0;
 sq2_trigger[80] = 0;
 sq2_trigger[81] = 0;
 sq2_trigger[82] = 0;
 sq2_trigger[83] = 0;
 sq2_trigger[84] = 1.0;
 sq2_trigger[85] = 0;
 sq2_trigger[86] = 0;
 sq2_trigger[87] = 0;
 sq2_trigger[88] = 1.0;
 sq2_trigger[89] = 0;
 sq2_trigger[90] = 0;
 sq2_trigger[91] = 0;
 sq2_trigger[92] = 1.0;
 sq2_trigger[93] = 0;
 sq2_trigger[94] = 0;
 sq2_trigger[95] = 0;
 sq2_trigger[96] = 1.0;
 sq2_trigger[97] = 0;
 sq2_trigger[98] = 0;
 sq2_trigger[99] = 0;
 sq2_trigger[100] = 0;
 sq2_trigger[101] = 0;
 sq2_trigger[102] = 1.0;
 sq2_trigger[103] = 0;
 sq2_trigger[104] = 0;
 sq2_trigger[105] = 0;
 sq2_trigger[106] = 0;
 sq2_trigger[107] = 0;
 sq2_trigger[108] = 1.0;
 sq2_trigger[109] = 0;
 sq2_trigger[110] = 0;
 sq2_trigger[111] = 1.0;
 sq2_trigger[112] = 0;
 sq2_trigger[113] = 0;
 sq2_trigger[114] = 1.0;
 sq2_trigger[115] = 0;
 sq2_trigger[116] = 0;
 sq2_trigger[117] = 1.0;
 sq2_trigger[118] = 0;
 sq2_trigger[119] = 0;
 sq2_trigger[120] = 1.0;
 sq2_trigger[121] = 0;
 sq2_trigger[122] = 0;
 sq2_trigger[123] = 0;
 sq2_trigger[124] = 1.0;
 sq2_trigger[125] = 0;
 sq2_trigger[126] = 0;
 sq2_trigger[127] = 0;
 sq2_trigger[128] = 1.0;
 sq2_trigger[129] = 0;
 sq2_trigger[130] = 0;
 sq2_trigger[131] = 0;
 sq2_trigger[132] = 1.0;
 sq2_trigger[133] = 0;
 sq2_trigger[134] = 0;
 sq2_trigger[135] = 0;
 sq2_trigger[136] = 1.0;
 sq2_trigger[137] = 0;
 sq2_trigger[138] = 0;
 sq2_trigger[139] = 0;
 sq2_trigger[140] = 1.0;
 sq2_trigger[141] = 0;
 sq2_trigger[142] = 0;
 sq2_trigger[143] = 0;
 sq2_trigger[144] = 1.0;
 sq2_trigger[145] = 0;
 sq2_trigger[146] = 0;
 sq2_trigger[147] = 0;
 sq2_trigger[148] = 0;
 sq2_trigger[149] = 0;
 sq2_trigger[150] = 0;
 sq2_trigger[151] = 0;
 sq2_trigger[152] = 1.0;
 sq2_trigger[153] = 0;
 sq2_trigger[154] = 0;
 sq2_trigger[155] = 0;
 sq2_trigger[156] = 1.0;
 sq2_trigger[157] = 0;
 sq2_trigger[158] = 0;
 sq2_trigger[159] = 0;
 sq2_trigger[160] = 1.0;
 sq2_trigger[161] = 0;
 sq2_trigger[162] = 0;
 sq2_trigger[163] = 0;
 sq2_trigger[164] = 1.0;
 sq2_trigger[165] = 0;
 sq2_trigger[166] = 0;
 sq2_trigger[167] = 0;
 sq2_trigger[168] = 1.0;
 sq2_trigger[169] = 0;
 sq2_trigger[170] = 0;
 sq2_trigger[171] = 0;
 sq2_trigger[172] = 0;
 sq2_trigger[173] = 0;
 sq2_trigger[174] = 0;
 sq2_trigger[175] = 0;
 sq2_trigger[176] = 1.0;
 sq2_trigger[177] = 0;
 sq2_trigger[178] = 0;
 sq2_trigger[179] = 0;
 sq2_trigger[180] = 1.0;
 sq2_trigger[181] = 0;
 sq2_trigger[182] = 0;
 sq2_trigger[183] = 0;
 sq2_trigger[184] = 1.0;
 sq2_trigger[185] = 0;
 sq2_trigger[186] = 0;
 sq2_trigger[187] = 0;
 sq2_trigger[188] = 1.0;
 sq2_trigger[189] = 0;
 sq2_trigger[190] = 0;
 sq2_trigger[191] = 0;
 sq2_trigger[192] = 1.0;
 sq2_trigger[193] = 0;
 sq2_trigger[194] = 0;
 sq2_trigger[195] = 0;
 sq2_trigger[196] = 0;
 sq2_trigger[197] = 0;
 sq2_trigger[198] = 1.0;
 sq2_trigger[199] = 0;
 sq2_trigger[200] = 0;
 sq2_trigger[201] = 1.0;
 sq2_trigger[202] = 0;
 sq2_trigger[203] = 0;
 sq2_trigger[204] = 1.0;
 sq2_trigger[205] = 0;
 sq2_trigger[206] = 0;
 sq2_trigger[207] = 0;
 sq2_trigger[208] = 0;
 sq2_trigger[209] = 0;
 sq2_trigger[210] = 1.0;
 sq2_trigger[211] = 0;
 sq2_trigger[212] = 0;
 sq2_trigger[213] = 1.0;
 sq2_trigger[214] = 0;
 sq2_trigger[215] = 0;
 sq2_trigger[216] = 1.0;
 sq2_trigger[217] = 0;
 sq2_trigger[218] = 0;
 sq2_trigger[219] = 0;
 sq2_trigger[220] = 0;
 sq2_trigger[221] = 0;
 sq2_trigger[222] = 0;
 sq2_trigger[223] = 0;
 sq2_trigger[224] = 0;
 sq2_trigger[225] = 0;
 sq2_trigger[226] = 0;
 sq2_trigger[227] = 0;
 sq2_trigger[228] = 1.0;
 sq2_trigger[229] = 0;
 sq2_trigger[230] = 0;
 sq2_trigger[231] = 0;
 sq2_trigger[232] = 0;
 sq2_trigger[233] = 0;
 sq2_trigger[234] = 1.0;
 sq2_trigger[235] = 0;
 sq2_trigger[236] = 0;
 sq2_trigger[237] = 0;
 sq2_trigger[238] = 0;
 sq2_trigger[239] = 0;
 sq2_trigger[240] = 1.0;
 sq2_trigger[241] = 0;
 sq2_trigger[242] = 0;
 sq2_trigger[243] = 0;
 sq2_trigger[244] = 0;
 sq2_trigger[245] = 0;
 sq2_trigger[246] = 1.0;
 sq2_trigger[247] = 0;
 sq2_trigger[248] = 0;
 sq2_trigger[249] = 1.0;
 sq2_trigger[250] = 0;
 sq2_trigger[251] = 0;
 sq2_trigger[252] = 1.0;
 sq2_trigger[253] = 0;
 sq2_trigger[254] = 0;
 sq2_trigger[255] = 0;
 sq2_trigger[256] = 0;
 sq2_trigger[257] = 0;
 sq2_trigger[258] = 1.0;
 sq2_trigger[259] = 0;
 sq2_trigger[260] = 0;
 sq2_trigger[261] = 1.0;
 sq2_trigger[262] = 0;
 sq2_trigger[263] = 0;
 sq2_trigger[264] = 1.0;
 sq2_trigger[265] = 0;
 sq2_trigger[266] = 0;
 sq2_trigger[267] = 0;
 sq2_trigger[268] = 0;
 sq2_trigger[269] = 0;
 sq2_trigger[270] = 0;
 sq2_trigger[271] = 0;
 sq2_trigger[272] = 0;
 sq2_trigger[273] = 0;
 sq2_trigger[274] = 0;
 sq2_trigger[275] = 0;
 sq2_trigger[276] = 1.0;
 sq2_trigger[277] = 0;
 sq2_trigger[278] = 0;
 sq2_trigger[279] = 0;
 sq2_trigger[280] = 0;
 sq2_trigger[281] = 0;
 sq2_trigger[282] = 1.0;
 sq2_trigger[283] = 0;
 sq2_trigger[284] = 0;
 sq2_trigger[285] = 0;
 sq2_trigger[286] = 0;
 sq2_trigger[287] = 0;
 sq2_trigger[288] = 1.0;
 sq2_trigger[289] = 0;
 sq2_trigger[290] = 0;
 sq2_trigger[291] = 0;
 sq2_trigger[292] = 0;
 sq2_trigger[293] = 0;
 sq2_trigger[294] = 0;
 sq2_trigger[295] = 0;
 sq2_trigger[296] = 0;
 sq2_trigger[297] = 0;
 sq2_trigger[298] = 0;
 sq2_trigger[299] = 0;
 sq2_trigger[300] = 1.0;
 sq2_trigger[301] = 0;
 sq2_trigger[302] = 0;
 sq2_trigger[303] = 0;
 sq2_trigger[304] = 0;
 sq2_trigger[305] = 0;
 sq2_trigger[306] = 1.0;
 sq2_trigger[307] = 0;
 sq2_trigger[308] = 0;
 sq2_trigger[309] = 1.0;
 sq2_trigger[310] = 0;
 sq2_trigger[311] = 0;
 sq2_trigger[312] = 1.0;
 sq2_trigger[313] = 0;
 sq2_trigger[314] = 0;
 sq2_trigger[315] = 0;
 sq2_trigger[316] = 0;
 sq2_trigger[317] = 0;
 sq2_trigger[318] = 1.0;
 sq2_trigger[319] = 0;
 sq2_trigger[320] = 0;
 sq2_trigger[321] = 1.0;
 sq2_trigger[322] = 0;
 sq2_trigger[323] = 0;
 sq2_trigger[324] = 1.0;
 sq2_trigger[325] = 0;
 sq2_trigger[326] = 0;
 sq2_trigger[327] = 0;
 sq2_trigger[328] = 0;
 sq2_trigger[329] = 0;
 sq2_trigger[330] = 1.0;
 sq2_trigger[331] = 0;
 sq2_trigger[332] = 0;
 sq2_trigger[333] = 0;
 sq2_trigger[334] = 0;
 sq2_trigger[335] = 0;
 sq2_trigger[336] = 1.0;
 sq2_trigger[337] = 0;
 sq2_trigger[338] = 0;
 sq2_trigger[339] = 0;
 sq2_trigger[340] = 0;
 sq2_trigger[341] = 0;
 sq2_trigger[342] = 0;
 sq2_trigger[343] = 0;
 sq2_trigger[344] = 0;
 sq2_trigger[345] = 0;
 sq2_trigger[346] = 0;
 sq2_trigger[347] = 0;
 sq2_trigger[348] = 0;
 sq2_trigger[349] = 0;
 sq2_trigger[350] = 0;
 sq2_trigger[351] = 0;
 sq2_trigger[352] = 0;
 sq2_trigger[353] = 0;
 sq2_trigger[354] = 0;
 sq2_trigger[355] = 0;
 sq2_trigger[356] = 0;
 sq2_trigger[357] = 0;
 sq2_trigger[358] = 0;
 sq2_trigger[359] = 0;
 sq2_trigger[360] = 0;
 sq2_trigger[361] = 0;
 sq2_trigger[362] = 0;
 sq2_trigger[363] = 0;
 sq2_trigger[364] = 0;
 sq2_trigger[365] = 0;
 sq2_trigger[366] = 0;
 sq2_trigger[367] = 0;
 sq2_trigger[368] = 0;
 sq2_trigger[369] = 0;
 sq2_trigger[370] = 0;
 sq2_trigger[371] = 0;
 sq2_trigger[372] = 0;
 sq2_trigger[373] = 0;
 sq2_trigger[374] = 0;
 sq2_trigger[375] = 0;
 sq2_trigger[376] = 0;
 sq2_trigger[377] = 0;
 sq2_trigger[378] = 0;
 sq2_lenEnable[0] = 1.0;
 sq2_lenEnable[1] = 1.0;
 sq2_lenEnable[2] = 1.0;
 sq2_lenEnable[3] = 1.0;
 sq2_lenEnable[4] = 1.0;
 sq2_lenEnable[5] = 1.0;
 sq2_lenEnable[6] = 1.0;
 sq2_lenEnable[7] = 1.0;
 sq2_lenEnable[8] = 1.0;
 sq2_lenEnable[9] = 1.0;
 sq2_lenEnable[10] = 1.0;
 sq2_lenEnable[11] = 1.0;
 sq2_lenEnable[12] = 1.0;
 sq2_lenEnable[13] = 1.0;
 sq2_lenEnable[14] = 1.0;
 sq2_lenEnable[15] = 1.0;
 sq2_lenEnable[16] = 1.0;
 sq2_lenEnable[17] = 1.0;
 sq2_lenEnable[18] = 1.0;
 sq2_lenEnable[19] = 1.0;
 sq2_lenEnable[20] = 1.0;
 sq2_lenEnable[21] = 1.0;
 sq2_lenEnable[22] = 1.0;
 sq2_lenEnable[23] = 1.0;
 sq2_lenEnable[24] = 1.0;
 sq2_lenEnable[25] = 1.0;
 sq2_lenEnable[26] = 1.0;
 sq2_lenEnable[27] = 1.0;
 sq2_lenEnable[28] = 1.0;
 sq2_lenEnable[29] = 1.0;
 sq2_lenEnable[30] = 1.0;
 sq2_lenEnable[31] = 1.0;
 sq2_lenEnable[32] = 1.0;
 sq2_lenEnable[33] = 1.0;
 sq2_lenEnable[34] = 1.0;
 sq2_lenEnable[35] = 1.0;
 sq2_lenEnable[36] = 1.0;
 sq2_lenEnable[37] = 1.0;
 sq2_lenEnable[38] = 1.0;
 sq2_lenEnable[39] = 1.0;
 sq2_lenEnable[40] = 1.0;
 sq2_lenEnable[41] = 1.0;
 sq2_lenEnable[42] = 1.0;
 sq2_lenEnable[43] = 1.0;
 sq2_lenEnable[44] = 1.0;
 sq2_lenEnable[45] = 1.0;
 sq2_lenEnable[46] = 1.0;
 sq2_lenEnable[47] = 1.0;
 sq2_lenEnable[48] = 1.0;
 sq2_lenEnable[49] = 1.0;
 sq2_lenEnable[50] = 1.0;
 sq2_lenEnable[51] = 1.0;
 sq2_lenEnable[52] = 1.0;
 sq2_lenEnable[53] = 1.0;
 sq2_lenEnable[54] = 1.0;
 sq2_lenEnable[55] = 1.0;
 sq2_lenEnable[56] = 1.0;
 sq2_lenEnable[57] = 1.0;
 sq2_lenEnable[58] = 1.0;
 sq2_lenEnable[59] = 1.0;
 sq2_lenEnable[60] = 1.0;
 sq2_lenEnable[61] = 1.0;
 sq2_lenEnable[62] = 1.0;
 sq2_lenEnable[63] = 1.0;
 sq2_lenEnable[64] = 1.0;
 sq2_lenEnable[65] = 1.0;
 sq2_lenEnable[66] = 1.0;
 sq2_lenEnable[67] = 1.0;
 sq2_lenEnable[68] = 1.0;
 sq2_lenEnable[69] = 1.0;
 sq2_lenEnable[70] = 1.0;
 sq2_lenEnable[71] = 1.0;
 sq2_lenEnable[72] = 1.0;
 sq2_lenEnable[73] = 1.0;
 sq2_lenEnable[74] = 1.0;
 sq2_lenEnable[75] = 1.0;
 sq2_lenEnable[76] = 1.0;
 sq2_lenEnable[77] = 1.0;
 sq2_lenEnable[78] = 1.0;
 sq2_lenEnable[79] = 1.0;
 sq2_lenEnable[80] = 1.0;
 sq2_lenEnable[81] = 1.0;
 sq2_lenEnable[82] = 1.0;
 sq2_lenEnable[83] = 1.0;
 sq2_lenEnable[84] = 1.0;
 sq2_lenEnable[85] = 1.0;
 sq2_lenEnable[86] = 1.0;
 sq2_lenEnable[87] = 1.0;
 sq2_lenEnable[88] = 1.0;
 sq2_lenEnable[89] = 1.0;
 sq2_lenEnable[90] = 1.0;
 sq2_lenEnable[91] = 1.0;
 sq2_lenEnable[92] = 1.0;
 sq2_lenEnable[93] = 1.0;
 sq2_lenEnable[94] = 1.0;
 sq2_lenEnable[95] = 1.0;
 sq2_lenEnable[96] = 1.0;
 sq2_lenEnable[97] = 1.0;
 sq2_lenEnable[98] = 1.0;
 sq2_lenEnable[99] = 1.0;
 sq2_lenEnable[100] = 1.0;
 sq2_lenEnable[101] = 1.0;
 sq2_lenEnable[102] = 1.0;
 sq2_lenEnable[103] = 1.0;
 sq2_lenEnable[104] = 1.0;
 sq2_lenEnable[105] = 1.0;
 sq2_lenEnable[106] = 1.0;
 sq2_lenEnable[107] = 1.0;
 sq2_lenEnable[108] = 1.0;
 sq2_lenEnable[109] = 1.0;
 sq2_lenEnable[110] = 1.0;
 sq2_lenEnable[111] = 1.0;
 sq2_lenEnable[112] = 1.0;
 sq2_lenEnable[113] = 1.0;
 sq2_lenEnable[114] = 1.0;
 sq2_lenEnable[115] = 1.0;
 sq2_lenEnable[116] = 1.0;
 sq2_lenEnable[117] = 1.0;
 sq2_lenEnable[118] = 1.0;
 sq2_lenEnable[119] = 1.0;
 sq2_lenEnable[120] = 1.0;
 sq2_lenEnable[121] = 1.0;
 sq2_lenEnable[122] = 1.0;
 sq2_lenEnable[123] = 1.0;
 sq2_lenEnable[124] = 1.0;
 sq2_lenEnable[125] = 1.0;
 sq2_lenEnable[126] = 1.0;
 sq2_lenEnable[127] = 1.0;
 sq2_lenEnable[128] = 1.0;
 sq2_lenEnable[129] = 1.0;
 sq2_lenEnable[130] = 1.0;
 sq2_lenEnable[131] = 1.0;
 sq2_lenEnable[132] = 1.0;
 sq2_lenEnable[133] = 1.0;
 sq2_lenEnable[134] = 1.0;
 sq2_lenEnable[135] = 1.0;
 sq2_lenEnable[136] = 1.0;
 sq2_lenEnable[137] = 1.0;
 sq2_lenEnable[138] = 1.0;
 sq2_lenEnable[139] = 1.0;
 sq2_lenEnable[140] = 1.0;
 sq2_lenEnable[141] = 1.0;
 sq2_lenEnable[142] = 1.0;
 sq2_lenEnable[143] = 1.0;
 sq2_lenEnable[144] = 1.0;
 sq2_lenEnable[145] = 1.0;
 sq2_lenEnable[146] = 1.0;
 sq2_lenEnable[147] = 1.0;
 sq2_lenEnable[148] = 1.0;
 sq2_lenEnable[149] = 1.0;
 sq2_lenEnable[150] = 1.0;
 sq2_lenEnable[151] = 1.0;
 sq2_lenEnable[152] = 1.0;
 sq2_lenEnable[153] = 1.0;
 sq2_lenEnable[154] = 1.0;
 sq2_lenEnable[155] = 1.0;
 sq2_lenEnable[156] = 1.0;
 sq2_lenEnable[157] = 1.0;
 sq2_lenEnable[158] = 1.0;
 sq2_lenEnable[159] = 1.0;
 sq2_lenEnable[160] = 1.0;
 sq2_lenEnable[161] = 1.0;
 sq2_lenEnable[162] = 1.0;
 sq2_lenEnable[163] = 1.0;
 sq2_lenEnable[164] = 1.0;
 sq2_lenEnable[165] = 1.0;
 sq2_lenEnable[166] = 1.0;
 sq2_lenEnable[167] = 1.0;
 sq2_lenEnable[168] = 1.0;
 sq2_lenEnable[169] = 1.0;
 sq2_lenEnable[170] = 1.0;
 sq2_lenEnable[171] = 1.0;
 sq2_lenEnable[172] = 1.0;
 sq2_lenEnable[173] = 1.0;
 sq2_lenEnable[174] = 1.0;
 sq2_lenEnable[175] = 1.0;
 sq2_lenEnable[176] = 1.0;
 sq2_lenEnable[177] = 1.0;
 sq2_lenEnable[178] = 1.0;
 sq2_lenEnable[179] = 1.0;
 sq2_lenEnable[180] = 1.0;
 sq2_lenEnable[181] = 1.0;
 sq2_lenEnable[182] = 1.0;
 sq2_lenEnable[183] = 1.0;
 sq2_lenEnable[184] = 1.0;
 sq2_lenEnable[185] = 1.0;
 sq2_lenEnable[186] = 1.0;
 sq2_lenEnable[187] = 1.0;
 sq2_lenEnable[188] = 1.0;
 sq2_lenEnable[189] = 1.0;
 sq2_lenEnable[190] = 1.0;
 sq2_lenEnable[191] = 1.0;
 sq2_lenEnable[192] = 1.0;
 sq2_lenEnable[193] = 1.0;
 sq2_lenEnable[194] = 1.0;
 sq2_lenEnable[195] = 1.0;
 sq2_lenEnable[196] = 1.0;
 sq2_lenEnable[197] = 1.0;
 sq2_lenEnable[198] = 1.0;
 sq2_lenEnable[199] = 1.0;
 sq2_lenEnable[200] = 1.0;
 sq2_lenEnable[201] = 1.0;
 sq2_lenEnable[202] = 1.0;
 sq2_lenEnable[203] = 1.0;
 sq2_lenEnable[204] = 1.0;
 sq2_lenEnable[205] = 1.0;
 sq2_lenEnable[206] = 1.0;
 sq2_lenEnable[207] = 1.0;
 sq2_lenEnable[208] = 1.0;
 sq2_lenEnable[209] = 1.0;
 sq2_lenEnable[210] = 1.0;
 sq2_lenEnable[211] = 1.0;
 sq2_lenEnable[212] = 1.0;
 sq2_lenEnable[213] = 1.0;
 sq2_lenEnable[214] = 1.0;
 sq2_lenEnable[215] = 1.0;
 sq2_lenEnable[216] = 1.0;
 sq2_lenEnable[217] = 1.0;
 sq2_lenEnable[218] = 1.0;
 sq2_lenEnable[219] = 1.0;
 sq2_lenEnable[220] = 1.0;
 sq2_lenEnable[221] = 1.0;
 sq2_lenEnable[222] = 1.0;
 sq2_lenEnable[223] = 1.0;
 sq2_lenEnable[224] = 1.0;
 sq2_lenEnable[225] = 1.0;
 sq2_lenEnable[226] = 1.0;
 sq2_lenEnable[227] = 1.0;
 sq2_lenEnable[228] = 1.0;
 sq2_lenEnable[229] = 1.0;
 sq2_lenEnable[230] = 1.0;
 sq2_lenEnable[231] = 1.0;
 sq2_lenEnable[232] = 1.0;
 sq2_lenEnable[233] = 1.0;
 sq2_lenEnable[234] = 1.0;
 sq2_lenEnable[235] = 1.0;
 sq2_lenEnable[236] = 1.0;
 sq2_lenEnable[237] = 1.0;
 sq2_lenEnable[238] = 1.0;
 sq2_lenEnable[239] = 1.0;
 sq2_lenEnable[240] = 1.0;
 sq2_lenEnable[241] = 1.0;
 sq2_lenEnable[242] = 1.0;
 sq2_lenEnable[243] = 1.0;
 sq2_lenEnable[244] = 1.0;
 sq2_lenEnable[245] = 1.0;
 sq2_lenEnable[246] = 1.0;
 sq2_lenEnable[247] = 1.0;
 sq2_lenEnable[248] = 1.0;
 sq2_lenEnable[249] = 1.0;
 sq2_lenEnable[250] = 1.0;
 sq2_lenEnable[251] = 1.0;
 sq2_lenEnable[252] = 1.0;
 sq2_lenEnable[253] = 1.0;
 sq2_lenEnable[254] = 1.0;
 sq2_lenEnable[255] = 1.0;
 sq2_lenEnable[256] = 1.0;
 sq2_lenEnable[257] = 1.0;
 sq2_lenEnable[258] = 1.0;
 sq2_lenEnable[259] = 1.0;
 sq2_lenEnable[260] = 1.0;
 sq2_lenEnable[261] = 1.0;
 sq2_lenEnable[262] = 1.0;
 sq2_lenEnable[263] = 1.0;
 sq2_lenEnable[264] = 1.0;
 sq2_lenEnable[265] = 1.0;
 sq2_lenEnable[266] = 1.0;
 sq2_lenEnable[267] = 1.0;
 sq2_lenEnable[268] = 1.0;
 sq2_lenEnable[269] = 1.0;
 sq2_lenEnable[270] = 1.0;
 sq2_lenEnable[271] = 1.0;
 sq2_lenEnable[272] = 1.0;
 sq2_lenEnable[273] = 1.0;
 sq2_lenEnable[274] = 1.0;
 sq2_lenEnable[275] = 1.0;
 sq2_lenEnable[276] = 1.0;
 sq2_lenEnable[277] = 1.0;
 sq2_lenEnable[278] = 1.0;
 sq2_lenEnable[279] = 1.0;
 sq2_lenEnable[280] = 1.0;
 sq2_lenEnable[281] = 1.0;
 sq2_lenEnable[282] = 1.0;
 sq2_lenEnable[283] = 1.0;
 sq2_lenEnable[284] = 1.0;
 sq2_lenEnable[285] = 1.0;
 sq2_lenEnable[286] = 1.0;
 sq2_lenEnable[287] = 1.0;
 sq2_lenEnable[288] = 1.0;
 sq2_lenEnable[289] = 1.0;
 sq2_lenEnable[290] = 1.0;
 sq2_lenEnable[291] = 1.0;
 sq2_lenEnable[292] = 1.0;
 sq2_lenEnable[293] = 1.0;
 sq2_lenEnable[294] = 1.0;
 sq2_lenEnable[295] = 1.0;
 sq2_lenEnable[296] = 1.0;
 sq2_lenEnable[297] = 1.0;
 sq2_lenEnable[298] = 1.0;
 sq2_lenEnable[299] = 1.0;
 sq2_lenEnable[300] = 1.0;
 sq2_lenEnable[301] = 1.0;
 sq2_lenEnable[302] = 1.0;
 sq2_lenEnable[303] = 1.0;
 sq2_lenEnable[304] = 1.0;
 sq2_lenEnable[305] = 1.0;
 sq2_lenEnable[306] = 1.0;
 sq2_lenEnable[307] = 1.0;
 sq2_lenEnable[308] = 1.0;
 sq2_lenEnable[309] = 1.0;
 sq2_lenEnable[310] = 1.0;
 sq2_lenEnable[311] = 1.0;
 sq2_lenEnable[312] = 1.0;
 sq2_lenEnable[313] = 1.0;
 sq2_lenEnable[314] = 1.0;
 sq2_lenEnable[315] = 1.0;
 sq2_lenEnable[316] = 1.0;
 sq2_lenEnable[317] = 1.0;
 sq2_lenEnable[318] = 1.0;
 sq2_lenEnable[319] = 1.0;
 sq2_lenEnable[320] = 1.0;
 sq2_lenEnable[321] = 1.0;
 sq2_lenEnable[322] = 1.0;
 sq2_lenEnable[323] = 1.0;
 sq2_lenEnable[324] = 1.0;
 sq2_lenEnable[325] = 1.0;
 sq2_lenEnable[326] = 1.0;
 sq2_lenEnable[327] = 1.0;
 sq2_lenEnable[328] = 1.0;
 sq2_lenEnable[329] = 1.0;
 sq2_lenEnable[330] = 1.0;
 sq2_lenEnable[331] = 1.0;
 sq2_lenEnable[332] = 1.0;
 sq2_lenEnable[333] = 1.0;
 sq2_lenEnable[334] = 1.0;
 sq2_lenEnable[335] = 1.0;
 sq2_lenEnable[336] = 1.0;
 sq2_lenEnable[337] = 1.0;
 sq2_lenEnable[338] = 1.0;
 sq2_lenEnable[339] = 1.0;
 sq2_lenEnable[340] = 1.0;
 sq2_lenEnable[341] = 1.0;
 sq2_lenEnable[342] = 1.0;
 sq2_lenEnable[343] = 1.0;
 sq2_lenEnable[344] = 1.0;
 sq2_lenEnable[345] = 1.0;
 sq2_lenEnable[346] = 1.0;
 sq2_lenEnable[347] = 1.0;
 sq2_lenEnable[348] = 1.0;
 sq2_lenEnable[349] = 1.0;
 sq2_lenEnable[350] = 1.0;
 sq2_lenEnable[351] = 1.0;
 sq2_lenEnable[352] = 1.0;
 sq2_lenEnable[353] = 1.0;
 sq2_lenEnable[354] = 1.0;
 sq2_lenEnable[355] = 1.0;
 sq2_lenEnable[356] = 1.0;
 sq2_lenEnable[357] = 1.0;
 sq2_lenEnable[358] = 1.0;
 sq2_lenEnable[359] = 1.0;
 sq2_lenEnable[360] = 1.0;
 sq2_lenEnable[361] = 1.0;
 sq2_lenEnable[362] = 1.0;
 sq2_lenEnable[363] = 1.0;
 sq2_lenEnable[364] = 1.0;
 sq2_lenEnable[365] = 1.0;
 sq2_lenEnable[366] = 1.0;
 sq2_lenEnable[367] = 1.0;
 sq2_lenEnable[368] = 1.0;
 sq2_lenEnable[369] = 1.0;
 sq2_lenEnable[370] = 1.0;
 sq2_lenEnable[371] = 1.0;
 sq2_lenEnable[372] = 1.0;
 sq2_lenEnable[373] = 1.0;
 sq2_lenEnable[374] = 1.0;
 sq2_lenEnable[375] = 1.0;
 sq2_lenEnable[376] = 1.0;
 sq2_lenEnable[377] = 1.0;
 sq2_lenEnable[378] = 1.0;


	end

endmodule
