`include "pulseChannel1.v"
`include "swDac.v"

`define PERIOD 4194304/16
`define LENGTH 10'd1023
`define PLAYBACK_LENGTH 10'd10
`define LONGREG reg [`LENGTH:0]

module gameboy();


	reg [31:0] [3:0] waveTable;

	// Square 1
	`LONGREG [2:0] sq1_swpPd;
	`LONGREG sq1_negate;
	`LONGREG [2:0] sq1_shift;
	`LONGREG [1:0] sq1_duty;
	`LONGREG [5:0] sq1_lenLoad;
	`LONGREG [3:0] sq1_startVol;
	`LONGREG sq1_envAdd;
	`LONGREG [2:0] sq1_period;
	`LONGREG [10:0] sq1_freq;
	`LONGREG sq1_trigger;
	`LONGREG sq1_lenEnable;

	wire clk; baseClk baseclk(clk);
	wire clk256; fixedTimer #(16384) tmr256(clk, clk256);
	wire clk128; fixedTimer #(2) tmr128(clk256, clk128);
	wire clk64; fixedTimer #(2) tmr64(clk128, clk64);

	wire clkT; fixedTimer #(`PERIOD) tmrT(clk, clkT);
	reg [$clog2(`LENGTH)-1:0] t;
	always @(posedge clkT) begin
		if (t < `PLAYBACK_LENGTH) t += 1;
		else $finish;
	end

	wire [3:0] sq1_out;
	pulseChannel1 pc1(clk, clk256, clk128, clk64, sq1_swpPd[t], sq1_negate[t], sq1_shift[t], sq1_freq[t], sq1_lenLoad[t], sq1_duty[t], sq1_startVol[t], sq1_period[t], sq1_trigger[t], sq1_lenEnable[t], sq1_envAdd[t], sq1_out);

	reg [4:0] ii; // Fill in the wave table with a triangle wave

	swDac dac(sq1_out, sq1_out);

	initial begin
		t = 0;

		for (ii = 0; ii < 16; ii++) waveTable[ii] = {ii[3:0]};
		for (ii = 0; ii < 16; ii++) waveTable[ii+5'd16] = 4'd0 - {ii[3:0]};

sq1_swpPd[0] <= 0.0; sq1_swpPd[1] <= 0.0; sq1_swpPd[2] <= 0.0; sq1_swpPd[3] <= 0.0; sq1_swpPd[4] <= 0.0; sq1_swpPd[5] <= 0.0; sq1_swpPd[6] <= 0.0; sq1_swpPd[7] <= 0.0; sq1_swpPd[8] <= 0.0; sq1_swpPd[9] <= 0.0; sq1_swpPd[10] <= 0.0; sq1_swpPd[11] <= 0.0; sq1_swpPd[12] <= 0.0; sq1_swpPd[13] <= 0.0; sq1_swpPd[14] <= 0.0; sq1_swpPd[15] <= 0.0; sq1_swpPd[16] <= 0.0; sq1_swpPd[17] <= 0.0; sq1_swpPd[18] <= 0.0; sq1_swpPd[19] <= 0.0; sq1_swpPd[20] <= 0.0; sq1_swpPd[21] <= 0.0; sq1_swpPd[22] <= 0.0; sq1_swpPd[23] <= 0.0; sq1_swpPd[24] <= 0.0; sq1_swpPd[25] <= 0.0; sq1_swpPd[26] <= 0.0; sq1_swpPd[27] <= 0.0; sq1_swpPd[28] <= 0.0; sq1_swpPd[29] <= 0.0; sq1_swpPd[30] <= 0.0; sq1_swpPd[31] <= 0.0; sq1_swpPd[32] <= 0.0; sq1_swpPd[33] <= 0.0; sq1_swpPd[34] <= 0.0; sq1_swpPd[35] <= 0.0; sq1_swpPd[36] <= 0.0; sq1_swpPd[37] <= 0.0; sq1_swpPd[38] <= 0.0; sq1_swpPd[39] <= 0.0; sq1_swpPd[40] <= 0.0; sq1_swpPd[41] <= 0.0; sq1_swpPd[42] <= 0.0; sq1_swpPd[43] <= 0.0; sq1_swpPd[44] <= 0.0; sq1_swpPd[45] <= 0.0; sq1_swpPd[46] <= 0.0; sq1_swpPd[47] <= 0.0; sq1_swpPd[48] <= 0.0; sq1_swpPd[49] <= 0.0; sq1_swpPd[50] <= 0.0; sq1_swpPd[51] <= 0.0; sq1_swpPd[52] <= 0.0; sq1_swpPd[53] <= 0.0; sq1_swpPd[54] <= 0.0; sq1_swpPd[55] <= 0.0; sq1_swpPd[56] <= 0.0; sq1_swpPd[57] <= 0.0; sq1_swpPd[58] <= 0.0; sq1_swpPd[59] <= 0.0; sq1_swpPd[60] <= 0.0; sq1_swpPd[61] <= 0.0; sq1_swpPd[62] <= 0.0; sq1_swpPd[63] <= 0.0; sq1_swpPd[64] <= 0.0; sq1_swpPd[65] <= 0.0; sq1_swpPd[66] <= 0.0; sq1_swpPd[67] <= 0.0; sq1_swpPd[68] <= 0.0; sq1_swpPd[69] <= 0.0; sq1_swpPd[70] <= 0.0; sq1_swpPd[71] <= 0.0; sq1_swpPd[72] <= 0.0; sq1_swpPd[73] <= 0.0; sq1_swpPd[74] <= 0.0; sq1_swpPd[75] <= 0.0; sq1_swpPd[76] <= 0.0; sq1_swpPd[77] <= 0.0; sq1_swpPd[78] <= 0.0; sq1_swpPd[79] <= 0.0; sq1_swpPd[80] <= 0.0; sq1_swpPd[81] <= 0.0; sq1_swpPd[82] <= 0.0; sq1_swpPd[83] <= 0.0; sq1_swpPd[84] <= 0.0; sq1_swpPd[85] <= 0.0; sq1_swpPd[86] <= 0.0; sq1_swpPd[87] <= 0.0; sq1_swpPd[88] <= 0.0; sq1_swpPd[89] <= 0.0; sq1_swpPd[90] <= 0.0; sq1_swpPd[91] <= 0.0; sq1_swpPd[92] <= 0.0; sq1_swpPd[93] <= 0.0; sq1_swpPd[94] <= 0.0; sq1_swpPd[95] <= 0.0; sq1_swpPd[96] <= 0.0; sq1_swpPd[97] <= 0.0; sq1_swpPd[98] <= 0.0; sq1_swpPd[99] <= 0.0; sq1_swpPd[100] <= 0.0; sq1_swpPd[101] <= 0.0; sq1_swpPd[102] <= 0.0; sq1_swpPd[103] <= 0.0; sq1_swpPd[104] <= 0.0; sq1_swpPd[105] <= 0.0; sq1_swpPd[106] <= 0.0; sq1_swpPd[107] <= 0.0; sq1_swpPd[108] <= 0.0; sq1_swpPd[109] <= 0.0; sq1_swpPd[110] <= 0.0; sq1_swpPd[111] <= 0.0; sq1_swpPd[112] <= 0.0; sq1_swpPd[113] <= 0.0; sq1_swpPd[114] <= 0.0; sq1_swpPd[115] <= 0.0; sq1_swpPd[116] <= 0.0; sq1_swpPd[117] <= 0.0; sq1_swpPd[118] <= 0.0; sq1_swpPd[119] <= 0.0; sq1_swpPd[120] <= 0.0; sq1_swpPd[121] <= 0.0; sq1_swpPd[122] <= 0.0; sq1_swpPd[123] <= 0.0; sq1_swpPd[124] <= 0.0; sq1_swpPd[125] <= 0.0; sq1_swpPd[126] <= 0.0; sq1_swpPd[127] <= 0.0; sq1_swpPd[128] <= 0.0; sq1_swpPd[129] <= 0.0; sq1_swpPd[130] <= 0.0; sq1_swpPd[131] <= 0.0; sq1_swpPd[132] <= 0.0; sq1_swpPd[133] <= 0.0; sq1_swpPd[134] <= 0.0; sq1_swpPd[135] <= 0.0; sq1_swpPd[136] <= 0.0; sq1_swpPd[137] <= 0.0; sq1_swpPd[138] <= 0.0; sq1_swpPd[139] <= 0.0; sq1_swpPd[140] <= 0.0; sq1_swpPd[141] <= 0.0; sq1_swpPd[142] <= 0.0; sq1_swpPd[143] <= 0.0; sq1_swpPd[144] <= 0.0; sq1_swpPd[145] <= 0.0; sq1_swpPd[146] <= 0.0; sq1_swpPd[147] <= 0.0; sq1_swpPd[148] <= 0.0; sq1_swpPd[149] <= 0.0; sq1_swpPd[150] <= 0.0; sq1_swpPd[151] <= 0.0; sq1_swpPd[152] <= 0.0; sq1_swpPd[153] <= 0.0; sq1_swpPd[154] <= 0.0; sq1_swpPd[155] <= 0.0; sq1_swpPd[156] <= 0.0; sq1_swpPd[157] <= 0.0; sq1_swpPd[158] <= 0.0; sq1_swpPd[159] <= 0.0; sq1_swpPd[160] <= 0.0; sq1_swpPd[161] <= 0.0; sq1_swpPd[162] <= 0.0; sq1_swpPd[163] <= 0.0; sq1_swpPd[164] <= 0.0; sq1_swpPd[165] <= 0.0; sq1_swpPd[166] <= 0.0; sq1_swpPd[167] <= 0.0; sq1_swpPd[168] <= 0.0; sq1_swpPd[169] <= 0.0; sq1_swpPd[170] <= 0.0; sq1_swpPd[171] <= 0.0; sq1_swpPd[172] <= 0.0; sq1_swpPd[173] <= 0.0; sq1_swpPd[174] <= 0.0; sq1_swpPd[175] <= 0.0; sq1_swpPd[176] <= 0.0; sq1_swpPd[177] <= 0.0; sq1_swpPd[178] <= 0.0; sq1_swpPd[179] <= 0.0; sq1_swpPd[180] <= 0.0; sq1_swpPd[181] <= 0.0; sq1_swpPd[182] <= 0.0; sq1_swpPd[183] <= 0.0; sq1_swpPd[184] <= 0.0; sq1_swpPd[185] <= 0.0; sq1_swpPd[186] <= 0.0; sq1_swpPd[187] <= 0.0; sq1_negate[0] <= 0.0; sq1_negate[1] <= 0.0; sq1_negate[2] <= 0.0; sq1_negate[3] <= 0.0; sq1_negate[4] <= 0.0; sq1_negate[5] <= 0.0; sq1_negate[6] <= 0.0; sq1_negate[7] <= 0.0; sq1_negate[8] <= 0.0; sq1_negate[9] <= 0.0; sq1_negate[10] <= 0.0; sq1_negate[11] <= 0.0; sq1_negate[12] <= 0.0; sq1_negate[13] <= 0.0; sq1_negate[14] <= 0.0; sq1_negate[15] <= 0.0; sq1_negate[16] <= 0.0; sq1_negate[17] <= 0.0; sq1_negate[18] <= 0.0; sq1_negate[19] <= 0.0; sq1_negate[20] <= 0.0; sq1_negate[21] <= 0.0; sq1_negate[22] <= 0.0; sq1_negate[23] <= 0.0; sq1_negate[24] <= 0.0; sq1_negate[25] <= 0.0; sq1_negate[26] <= 0.0; sq1_negate[27] <= 0.0; sq1_negate[28] <= 0.0; sq1_negate[29] <= 0.0; sq1_negate[30] <= 0.0; sq1_negate[31] <= 0.0; sq1_negate[32] <= 0.0; sq1_negate[33] <= 0.0; sq1_negate[34] <= 0.0; sq1_negate[35] <= 0.0; sq1_negate[36] <= 0.0; sq1_negate[37] <= 0.0; sq1_negate[38] <= 0.0; sq1_negate[39] <= 0.0; sq1_negate[40] <= 0.0; sq1_negate[41] <= 0.0; sq1_negate[42] <= 0.0; sq1_negate[43] <= 0.0; sq1_negate[44] <= 0.0; sq1_negate[45] <= 0.0; sq1_negate[46] <= 0.0; sq1_negate[47] <= 0.0; sq1_negate[48] <= 0.0; sq1_negate[49] <= 0.0; sq1_negate[50] <= 0.0; sq1_negate[51] <= 0.0; sq1_negate[52] <= 0.0; sq1_negate[53] <= 0.0; sq1_negate[54] <= 0.0; sq1_negate[55] <= 0.0; sq1_negate[56] <= 0.0; sq1_negate[57] <= 0.0; sq1_negate[58] <= 0.0; sq1_negate[59] <= 0.0; sq1_negate[60] <= 0.0; sq1_negate[61] <= 0.0; sq1_negate[62] <= 0.0; sq1_negate[63] <= 0.0; sq1_negate[64] <= 0.0; sq1_negate[65] <= 0.0; sq1_negate[66] <= 0.0; sq1_negate[67] <= 0.0; sq1_negate[68] <= 0.0; sq1_negate[69] <= 0.0; sq1_negate[70] <= 0.0; sq1_negate[71] <= 0.0; sq1_negate[72] <= 0.0; sq1_negate[73] <= 0.0; sq1_negate[74] <= 0.0; sq1_negate[75] <= 0.0; sq1_negate[76] <= 0.0; sq1_negate[77] <= 0.0; sq1_negate[78] <= 0.0; sq1_negate[79] <= 0.0; sq1_negate[80] <= 0.0; sq1_negate[81] <= 0.0; sq1_negate[82] <= 0.0; sq1_negate[83] <= 0.0; sq1_negate[84] <= 0.0; sq1_negate[85] <= 0.0; sq1_negate[86] <= 0.0; sq1_negate[87] <= 0.0; sq1_negate[88] <= 0.0; sq1_negate[89] <= 0.0; sq1_negate[90] <= 0.0; sq1_negate[91] <= 0.0; sq1_negate[92] <= 0.0; sq1_negate[93] <= 0.0; sq1_negate[94] <= 0.0; sq1_negate[95] <= 0.0; sq1_negate[96] <= 0.0; sq1_negate[97] <= 0.0; sq1_negate[98] <= 0.0; sq1_negate[99] <= 0.0; sq1_negate[100] <= 0.0; sq1_negate[101] <= 0.0; sq1_negate[102] <= 0.0; sq1_negate[103] <= 0.0; sq1_negate[104] <= 0.0; sq1_negate[105] <= 0.0; sq1_negate[106] <= 0.0; sq1_negate[107] <= 0.0; sq1_negate[108] <= 0.0; sq1_negate[109] <= 0.0; sq1_negate[110] <= 0.0; sq1_negate[111] <= 0.0; sq1_negate[112] <= 0.0; sq1_negate[113] <= 0.0; sq1_negate[114] <= 0.0; sq1_negate[115] <= 0.0; sq1_negate[116] <= 0.0; sq1_negate[117] <= 0.0; sq1_negate[118] <= 0.0; sq1_negate[119] <= 0.0; sq1_negate[120] <= 0.0; sq1_negate[121] <= 0.0; sq1_negate[122] <= 0.0; sq1_negate[123] <= 0.0; sq1_negate[124] <= 0.0; sq1_negate[125] <= 0.0; sq1_negate[126] <= 0.0; sq1_negate[127] <= 0.0; sq1_negate[128] <= 0.0; sq1_negate[129] <= 0.0; sq1_negate[130] <= 0.0; sq1_negate[131] <= 0.0; sq1_negate[132] <= 0.0; sq1_negate[133] <= 0.0; sq1_negate[134] <= 0.0; sq1_negate[135] <= 0.0; sq1_negate[136] <= 0.0; sq1_negate[137] <= 0.0; sq1_negate[138] <= 0.0; sq1_negate[139] <= 0.0; sq1_negate[140] <= 0.0; sq1_negate[141] <= 0.0; sq1_negate[142] <= 0.0; sq1_negate[143] <= 0.0; sq1_negate[144] <= 0.0; sq1_negate[145] <= 0.0; sq1_negate[146] <= 0.0; sq1_negate[147] <= 0.0; sq1_negate[148] <= 0.0; sq1_negate[149] <= 0.0; sq1_negate[150] <= 0.0; sq1_negate[151] <= 0.0; sq1_negate[152] <= 0.0; sq1_negate[153] <= 0.0; sq1_negate[154] <= 0.0; sq1_negate[155] <= 0.0; sq1_negate[156] <= 0.0; sq1_negate[157] <= 0.0; sq1_negate[158] <= 0.0; sq1_negate[159] <= 0.0; sq1_negate[160] <= 0.0; sq1_negate[161] <= 0.0; sq1_negate[162] <= 0.0; sq1_negate[163] <= 0.0; sq1_negate[164] <= 0.0; sq1_negate[165] <= 0.0; sq1_negate[166] <= 0.0; sq1_negate[167] <= 0.0; sq1_negate[168] <= 0.0; sq1_negate[169] <= 0.0; sq1_negate[170] <= 0.0; sq1_negate[171] <= 0.0; sq1_negate[172] <= 0.0; sq1_negate[173] <= 0.0; sq1_negate[174] <= 0.0; sq1_negate[175] <= 0.0; sq1_negate[176] <= 0.0; sq1_negate[177] <= 0.0; sq1_negate[178] <= 0.0; sq1_negate[179] <= 0.0; sq1_negate[180] <= 0.0; sq1_negate[181] <= 0.0; sq1_negate[182] <= 0.0; sq1_negate[183] <= 0.0; sq1_negate[184] <= 0.0; sq1_negate[185] <= 0.0; sq1_negate[186] <= 0.0; sq1_negate[187] <= 0.0; sq1_shift[0] <= 0.0; sq1_shift[1] <= 0.0; sq1_shift[2] <= 0.0; sq1_shift[3] <= 0.0; sq1_shift[4] <= 0.0; sq1_shift[5] <= 0.0; sq1_shift[6] <= 0.0; sq1_shift[7] <= 0.0; sq1_shift[8] <= 0.0; sq1_shift[9] <= 0.0; sq1_shift[10] <= 0.0; sq1_shift[11] <= 0.0; sq1_shift[12] <= 0.0; sq1_shift[13] <= 0.0; sq1_shift[14] <= 0.0; sq1_shift[15] <= 0.0; sq1_shift[16] <= 0.0; sq1_shift[17] <= 0.0; sq1_shift[18] <= 0.0; sq1_shift[19] <= 0.0; sq1_shift[20] <= 0.0; sq1_shift[21] <= 0.0; sq1_shift[22] <= 0.0; sq1_shift[23] <= 0.0; sq1_shift[24] <= 0.0; sq1_shift[25] <= 0.0; sq1_shift[26] <= 0.0; sq1_shift[27] <= 0.0; sq1_shift[28] <= 0.0; sq1_shift[29] <= 0.0; sq1_shift[30] <= 0.0; sq1_shift[31] <= 0.0; sq1_shift[32] <= 0.0; sq1_shift[33] <= 0.0; sq1_shift[34] <= 0.0; sq1_shift[35] <= 0.0; sq1_shift[36] <= 0.0; sq1_shift[37] <= 0.0; sq1_shift[38] <= 0.0; sq1_shift[39] <= 0.0; sq1_shift[40] <= 0.0; sq1_shift[41] <= 0.0; sq1_shift[42] <= 0.0; sq1_shift[43] <= 0.0; sq1_shift[44] <= 0.0; sq1_shift[45] <= 0.0; sq1_shift[46] <= 0.0; sq1_shift[47] <= 0.0; sq1_shift[48] <= 0.0; sq1_shift[49] <= 0.0; sq1_shift[50] <= 0.0; sq1_shift[51] <= 0.0; sq1_shift[52] <= 0.0; sq1_shift[53] <= 0.0; sq1_shift[54] <= 0.0; sq1_shift[55] <= 0.0; sq1_shift[56] <= 0.0; sq1_shift[57] <= 0.0; sq1_shift[58] <= 0.0; sq1_shift[59] <= 0.0; sq1_shift[60] <= 0.0; sq1_shift[61] <= 0.0; sq1_shift[62] <= 0.0; sq1_shift[63] <= 0.0; sq1_shift[64] <= 0.0; sq1_shift[65] <= 0.0; sq1_shift[66] <= 0.0; sq1_shift[67] <= 0.0; sq1_shift[68] <= 0.0; sq1_shift[69] <= 0.0; sq1_shift[70] <= 0.0; sq1_shift[71] <= 0.0; sq1_shift[72] <= 0.0; sq1_shift[73] <= 0.0; sq1_shift[74] <= 0.0; sq1_shift[75] <= 0.0; sq1_shift[76] <= 0.0; sq1_shift[77] <= 0.0; sq1_shift[78] <= 0.0; sq1_shift[79] <= 0.0; sq1_shift[80] <= 0.0; sq1_shift[81] <= 0.0; sq1_shift[82] <= 0.0; sq1_shift[83] <= 0.0; sq1_shift[84] <= 0.0; sq1_shift[85] <= 0.0; sq1_shift[86] <= 0.0; sq1_shift[87] <= 0.0; sq1_shift[88] <= 0.0; sq1_shift[89] <= 0.0; sq1_shift[90] <= 0.0; sq1_shift[91] <= 0.0; sq1_shift[92] <= 0.0; sq1_shift[93] <= 0.0; sq1_shift[94] <= 0.0; sq1_shift[95] <= 0.0; sq1_shift[96] <= 0.0; sq1_shift[97] <= 0.0; sq1_shift[98] <= 0.0; sq1_shift[99] <= 0.0; sq1_shift[100] <= 0.0; sq1_shift[101] <= 0.0; sq1_shift[102] <= 0.0; sq1_shift[103] <= 0.0; sq1_shift[104] <= 0.0; sq1_shift[105] <= 0.0; sq1_shift[106] <= 0.0; sq1_shift[107] <= 0.0; sq1_shift[108] <= 0.0; sq1_shift[109] <= 0.0; sq1_shift[110] <= 0.0; sq1_shift[111] <= 0.0; sq1_shift[112] <= 0.0; sq1_shift[113] <= 0.0; sq1_shift[114] <= 0.0; sq1_shift[115] <= 0.0; sq1_shift[116] <= 0.0; sq1_shift[117] <= 0.0; sq1_shift[118] <= 0.0; sq1_shift[119] <= 0.0; sq1_shift[120] <= 0.0; sq1_shift[121] <= 0.0; sq1_shift[122] <= 0.0; sq1_shift[123] <= 0.0; sq1_shift[124] <= 0.0; sq1_shift[125] <= 0.0; sq1_shift[126] <= 0.0; sq1_shift[127] <= 0.0; sq1_shift[128] <= 0.0; sq1_shift[129] <= 0.0; sq1_shift[130] <= 0.0; sq1_shift[131] <= 0.0; sq1_shift[132] <= 0.0; sq1_shift[133] <= 0.0; sq1_shift[134] <= 0.0; sq1_shift[135] <= 0.0; sq1_shift[136] <= 0.0; sq1_shift[137] <= 0.0; sq1_shift[138] <= 0.0; sq1_shift[139] <= 0.0; sq1_shift[140] <= 0.0; sq1_shift[141] <= 0.0; sq1_shift[142] <= 0.0; sq1_shift[143] <= 0.0; sq1_shift[144] <= 0.0; sq1_shift[145] <= 0.0; sq1_shift[146] <= 0.0; sq1_shift[147] <= 0.0; sq1_shift[148] <= 0.0; sq1_shift[149] <= 0.0; sq1_shift[150] <= 0.0; sq1_shift[151] <= 0.0; sq1_shift[152] <= 0.0; sq1_shift[153] <= 0.0; sq1_shift[154] <= 0.0; sq1_shift[155] <= 0.0; sq1_shift[156] <= 0.0; sq1_shift[157] <= 0.0; sq1_shift[158] <= 0.0; sq1_shift[159] <= 0.0; sq1_shift[160] <= 0.0; sq1_shift[161] <= 0.0; sq1_shift[162] <= 0.0; sq1_shift[163] <= 0.0; sq1_shift[164] <= 0.0; sq1_shift[165] <= 0.0; sq1_shift[166] <= 0.0; sq1_shift[167] <= 0.0; sq1_shift[168] <= 0.0; sq1_shift[169] <= 0.0; sq1_shift[170] <= 0.0; sq1_shift[171] <= 0.0; sq1_shift[172] <= 0.0; sq1_shift[173] <= 0.0; sq1_shift[174] <= 0.0; sq1_shift[175] <= 0.0; sq1_shift[176] <= 0.0; sq1_shift[177] <= 0.0; sq1_shift[178] <= 0.0; sq1_shift[179] <= 0.0; sq1_shift[180] <= 0.0; sq1_shift[181] <= 0.0; sq1_shift[182] <= 0.0; sq1_shift[183] <= 0.0; sq1_shift[184] <= 0.0; sq1_shift[185] <= 0.0; sq1_shift[186] <= 0.0; sq1_shift[187] <= 0.0; sq1_duty[0] <= 2.0; sq1_duty[1] <= 2.0; sq1_duty[2] <= 2.0; sq1_duty[3] <= 2.0; sq1_duty[4] <= 2.0; sq1_duty[5] <= 2.0; sq1_duty[6] <= 2.0; sq1_duty[7] <= 2.0; sq1_duty[8] <= 2.0; sq1_duty[9] <= 2.0; sq1_duty[10] <= 2.0; sq1_duty[11] <= 2.0; sq1_duty[12] <= 2.0; sq1_duty[13] <= 2.0; sq1_duty[14] <= 2.0; sq1_duty[15] <= 2.0; sq1_duty[16] <= 2.0; sq1_duty[17] <= 2.0; sq1_duty[18] <= 2.0; sq1_duty[19] <= 2.0; sq1_duty[20] <= 2.0; sq1_duty[21] <= 2.0; sq1_duty[22] <= 2.0; sq1_duty[23] <= 2.0; sq1_duty[24] <= 2.0; sq1_duty[25] <= 2.0; sq1_duty[26] <= 2.0; sq1_duty[27] <= 2.0; sq1_duty[28] <= 2.0; sq1_duty[29] <= 2.0; sq1_duty[30] <= 2.0; sq1_duty[31] <= 2.0; sq1_duty[32] <= 2.0; sq1_duty[33] <= 2.0; sq1_duty[34] <= 2.0; sq1_duty[35] <= 2.0; sq1_duty[36] <= 2.0; sq1_duty[37] <= 2.0; sq1_duty[38] <= 2.0; sq1_duty[39] <= 2.0; sq1_duty[40] <= 2.0; sq1_duty[41] <= 2.0; sq1_duty[42] <= 2.0; sq1_duty[43] <= 2.0; sq1_duty[44] <= 2.0; sq1_duty[45] <= 2.0; sq1_duty[46] <= 2.0; sq1_duty[47] <= 2.0; sq1_duty[48] <= 2.0; sq1_duty[49] <= 2.0; sq1_duty[50] <= 2.0; sq1_duty[51] <= 2.0; sq1_duty[52] <= 2.0; sq1_duty[53] <= 2.0; sq1_duty[54] <= 2.0; sq1_duty[55] <= 2.0; sq1_duty[56] <= 2.0; sq1_duty[57] <= 2.0; sq1_duty[58] <= 2.0; sq1_duty[59] <= 2.0; sq1_duty[60] <= 2.0; sq1_duty[61] <= 2.0; sq1_duty[62] <= 2.0; sq1_duty[63] <= 2.0; sq1_duty[64] <= 2.0; sq1_duty[65] <= 2.0; sq1_duty[66] <= 2.0; sq1_duty[67] <= 2.0; sq1_duty[68] <= 2.0; sq1_duty[69] <= 2.0; sq1_duty[70] <= 2.0; sq1_duty[71] <= 2.0; sq1_duty[72] <= 2.0; sq1_duty[73] <= 2.0; sq1_duty[74] <= 2.0; sq1_duty[75] <= 2.0; sq1_duty[76] <= 2.0; sq1_duty[77] <= 2.0; sq1_duty[78] <= 2.0; sq1_duty[79] <= 2.0; sq1_duty[80] <= 2.0; sq1_duty[81] <= 2.0; sq1_duty[82] <= 2.0; sq1_duty[83] <= 2.0; sq1_duty[84] <= 2.0; sq1_duty[85] <= 2.0; sq1_duty[86] <= 2.0; sq1_duty[87] <= 2.0; sq1_duty[88] <= 2.0; sq1_duty[89] <= 2.0; sq1_duty[90] <= 2.0; sq1_duty[91] <= 2.0; sq1_duty[92] <= 2.0; sq1_duty[93] <= 2.0; sq1_duty[94] <= 2.0; sq1_duty[95] <= 2.0; sq1_duty[96] <= 2.0; sq1_duty[97] <= 2.0; sq1_duty[98] <= 2.0; sq1_duty[99] <= 2.0; sq1_duty[100] <= 2.0; sq1_duty[101] <= 2.0; sq1_duty[102] <= 2.0; sq1_duty[103] <= 2.0; sq1_duty[104] <= 2.0; sq1_duty[105] <= 2.0; sq1_duty[106] <= 2.0; sq1_duty[107] <= 2.0; sq1_duty[108] <= 2.0; sq1_duty[109] <= 2.0; sq1_duty[110] <= 2.0; sq1_duty[111] <= 2.0; sq1_duty[112] <= 2.0; sq1_duty[113] <= 2.0; sq1_duty[114] <= 2.0; sq1_duty[115] <= 2.0; sq1_duty[116] <= 2.0; sq1_duty[117] <= 2.0; sq1_duty[118] <= 2.0; sq1_duty[119] <= 2.0; sq1_duty[120] <= 2.0; sq1_duty[121] <= 2.0; sq1_duty[122] <= 2.0; sq1_duty[123] <= 2.0; sq1_duty[124] <= 2.0; sq1_duty[125] <= 2.0; sq1_duty[126] <= 2.0; sq1_duty[127] <= 2.0; sq1_duty[128] <= 2.0; sq1_duty[129] <= 2.0; sq1_duty[130] <= 2.0; sq1_duty[131] <= 2.0; sq1_duty[132] <= 2.0; sq1_duty[133] <= 2.0; sq1_duty[134] <= 2.0; sq1_duty[135] <= 2.0; sq1_duty[136] <= 2.0; sq1_duty[137] <= 2.0; sq1_duty[138] <= 2.0; sq1_duty[139] <= 2.0; sq1_duty[140] <= 2.0; sq1_duty[141] <= 2.0; sq1_duty[142] <= 2.0; sq1_duty[143] <= 2.0; sq1_duty[144] <= 2.0; sq1_duty[145] <= 2.0; sq1_duty[146] <= 2.0; sq1_duty[147] <= 2.0; sq1_duty[148] <= 2.0; sq1_duty[149] <= 2.0; sq1_duty[150] <= 2.0; sq1_duty[151] <= 2.0; sq1_duty[152] <= 2.0; sq1_duty[153] <= 2.0; sq1_duty[154] <= 2.0; sq1_duty[155] <= 2.0; sq1_duty[156] <= 2.0; sq1_duty[157] <= 2.0; sq1_duty[158] <= 2.0; sq1_duty[159] <= 2.0; sq1_duty[160] <= 2.0; sq1_duty[161] <= 2.0; sq1_duty[162] <= 2.0; sq1_duty[163] <= 2.0; sq1_duty[164] <= 2.0; sq1_duty[165] <= 2.0; sq1_duty[166] <= 2.0; sq1_duty[167] <= 2.0; sq1_duty[168] <= 2.0; sq1_duty[169] <= 2.0; sq1_duty[170] <= 2.0; sq1_duty[171] <= 2.0; sq1_duty[172] <= 2.0; sq1_duty[173] <= 2.0; sq1_duty[174] <= 2.0; sq1_duty[175] <= 2.0; sq1_duty[176] <= 2.0; sq1_duty[177] <= 2.0; sq1_duty[178] <= 2.0; sq1_duty[179] <= 2.0; sq1_duty[180] <= 2.0; sq1_duty[181] <= 2.0; sq1_duty[182] <= 2.0; sq1_duty[183] <= 2.0; sq1_duty[184] <= 2.0; sq1_duty[185] <= 2.0; sq1_duty[186] <= 2.0; sq1_duty[187] <= 2.0; sq1_lenLoad[0] <= 32.0; sq1_lenLoad[1] <= 32.0; sq1_lenLoad[2] <= 32.0; sq1_lenLoad[3] <= 32.0; sq1_lenLoad[4] <= 32.0; sq1_lenLoad[5] <= 32.0; sq1_lenLoad[6] <= 32.0; sq1_lenLoad[7] <= 32.0; sq1_lenLoad[8] <= 32.0; sq1_lenLoad[9] <= 32.0; sq1_lenLoad[10] <= 32.0; sq1_lenLoad[11] <= 32.0; sq1_lenLoad[12] <= 32.0; sq1_lenLoad[13] <= 32.0; sq1_lenLoad[14] <= 32.0; sq1_lenLoad[15] <= 32.0; sq1_lenLoad[16] <= 32.0; sq1_lenLoad[17] <= 32.0; sq1_lenLoad[18] <= 32.0; sq1_lenLoad[19] <= 32.0; sq1_lenLoad[20] <= 32.0; sq1_lenLoad[21] <= 32.0; sq1_lenLoad[22] <= 32.0; sq1_lenLoad[23] <= 32.0; sq1_lenLoad[24] <= 32.0; sq1_lenLoad[25] <= 32.0; sq1_lenLoad[26] <= 32.0; sq1_lenLoad[27] <= 32.0; sq1_lenLoad[28] <= 32.0; sq1_lenLoad[29] <= 32.0; sq1_lenLoad[30] <= 32.0; sq1_lenLoad[31] <= 32.0; sq1_lenLoad[32] <= 32.0; sq1_lenLoad[33] <= 32.0; sq1_lenLoad[34] <= 32.0; sq1_lenLoad[35] <= 32.0; sq1_lenLoad[36] <= 32.0; sq1_lenLoad[37] <= 32.0; sq1_lenLoad[38] <= 32.0; sq1_lenLoad[39] <= 32.0; sq1_lenLoad[40] <= 32.0; sq1_lenLoad[41] <= 32.0; sq1_lenLoad[42] <= 32.0; sq1_lenLoad[43] <= 32.0; sq1_lenLoad[44] <= 32.0; sq1_lenLoad[45] <= 32.0; sq1_lenLoad[46] <= 32.0; sq1_lenLoad[47] <= 32.0; sq1_lenLoad[48] <= 32.0; sq1_lenLoad[49] <= 32.0; sq1_lenLoad[50] <= 32.0; sq1_lenLoad[51] <= 32.0; sq1_lenLoad[52] <= 32.0; sq1_lenLoad[53] <= 32.0; sq1_lenLoad[54] <= 32.0; sq1_lenLoad[55] <= 32.0; sq1_lenLoad[56] <= 32.0; sq1_lenLoad[57] <= 32.0; sq1_lenLoad[58] <= 32.0; sq1_lenLoad[59] <= 32.0; sq1_lenLoad[60] <= 32.0; sq1_lenLoad[61] <= 32.0; sq1_lenLoad[62] <= 32.0; sq1_lenLoad[63] <= 32.0; sq1_lenLoad[64] <= 32.0; sq1_lenLoad[65] <= 32.0; sq1_lenLoad[66] <= 32.0; sq1_lenLoad[67] <= 32.0; sq1_lenLoad[68] <= 32.0; sq1_lenLoad[69] <= 32.0; sq1_lenLoad[70] <= 32.0; sq1_lenLoad[71] <= 32.0; sq1_lenLoad[72] <= 32.0; sq1_lenLoad[73] <= 32.0; sq1_lenLoad[74] <= 32.0; sq1_lenLoad[75] <= 32.0; sq1_lenLoad[76] <= 32.0; sq1_lenLoad[77] <= 32.0; sq1_lenLoad[78] <= 32.0; sq1_lenLoad[79] <= 32.0; sq1_lenLoad[80] <= 32.0; sq1_lenLoad[81] <= 32.0; sq1_lenLoad[82] <= 32.0; sq1_lenLoad[83] <= 32.0; sq1_lenLoad[84] <= 32.0; sq1_lenLoad[85] <= 32.0; sq1_lenLoad[86] <= 32.0; sq1_lenLoad[87] <= 32.0; sq1_lenLoad[88] <= 32.0; sq1_lenLoad[89] <= 32.0; sq1_lenLoad[90] <= 32.0; sq1_lenLoad[91] <= 32.0; sq1_lenLoad[92] <= 32.0; sq1_lenLoad[93] <= 32.0; sq1_lenLoad[94] <= 32.0; sq1_lenLoad[95] <= 32.0; sq1_lenLoad[96] <= 32.0; sq1_lenLoad[97] <= 32.0; sq1_lenLoad[98] <= 32.0; sq1_lenLoad[99] <= 32.0; sq1_lenLoad[100] <= 32.0; sq1_lenLoad[101] <= 32.0; sq1_lenLoad[102] <= 32.0; sq1_lenLoad[103] <= 32.0; sq1_lenLoad[104] <= 32.0; sq1_lenLoad[105] <= 32.0; sq1_lenLoad[106] <= 32.0; sq1_lenLoad[107] <= 32.0; sq1_lenLoad[108] <= 32.0; sq1_lenLoad[109] <= 32.0; sq1_lenLoad[110] <= 32.0; sq1_lenLoad[111] <= 32.0; sq1_lenLoad[112] <= 32.0; sq1_lenLoad[113] <= 32.0; sq1_lenLoad[114] <= 32.0; sq1_lenLoad[115] <= 32.0; sq1_lenLoad[116] <= 32.0; sq1_lenLoad[117] <= 32.0; sq1_lenLoad[118] <= 32.0; sq1_lenLoad[119] <= 32.0; sq1_lenLoad[120] <= 32.0; sq1_lenLoad[121] <= 32.0; sq1_lenLoad[122] <= 32.0; sq1_lenLoad[123] <= 32.0; sq1_lenLoad[124] <= 32.0; sq1_lenLoad[125] <= 32.0; sq1_lenLoad[126] <= 32.0; sq1_lenLoad[127] <= 32.0; sq1_lenLoad[128] <= 32.0; sq1_lenLoad[129] <= 32.0; sq1_lenLoad[130] <= 32.0; sq1_lenLoad[131] <= 32.0; sq1_lenLoad[132] <= 32.0; sq1_lenLoad[133] <= 32.0; sq1_lenLoad[134] <= 32.0; sq1_lenLoad[135] <= 32.0; sq1_lenLoad[136] <= 32.0; sq1_lenLoad[137] <= 32.0; sq1_lenLoad[138] <= 32.0; sq1_lenLoad[139] <= 32.0; sq1_lenLoad[140] <= 32.0; sq1_lenLoad[141] <= 32.0; sq1_lenLoad[142] <= 32.0; sq1_lenLoad[143] <= 32.0; sq1_lenLoad[144] <= 32.0; sq1_lenLoad[145] <= 32.0; sq1_lenLoad[146] <= 32.0; sq1_lenLoad[147] <= 32.0; sq1_lenLoad[148] <= 32.0; sq1_lenLoad[149] <= 32.0; sq1_lenLoad[150] <= 32.0; sq1_lenLoad[151] <= 32.0; sq1_lenLoad[152] <= 32.0; sq1_lenLoad[153] <= 32.0; sq1_lenLoad[154] <= 32.0; sq1_lenLoad[155] <= 32.0; sq1_lenLoad[156] <= 32.0; sq1_lenLoad[157] <= 32.0; sq1_lenLoad[158] <= 32.0; sq1_lenLoad[159] <= 32.0; sq1_lenLoad[160] <= 32.0; sq1_lenLoad[161] <= 32.0; sq1_lenLoad[162] <= 32.0; sq1_lenLoad[163] <= 32.0; sq1_lenLoad[164] <= 32.0; sq1_lenLoad[165] <= 32.0; sq1_lenLoad[166] <= 32.0; sq1_lenLoad[167] <= 32.0; sq1_lenLoad[168] <= 32.0; sq1_lenLoad[169] <= 32.0; sq1_lenLoad[170] <= 32.0; sq1_lenLoad[171] <= 32.0; sq1_lenLoad[172] <= 32.0; sq1_lenLoad[173] <= 32.0; sq1_lenLoad[174] <= 32.0; sq1_lenLoad[175] <= 32.0; sq1_lenLoad[176] <= 32.0; sq1_lenLoad[177] <= 32.0; sq1_lenLoad[178] <= 32.0; sq1_lenLoad[179] <= 32.0; sq1_lenLoad[180] <= 32.0; sq1_lenLoad[181] <= 32.0; sq1_lenLoad[182] <= 32.0; sq1_lenLoad[183] <= 32.0; sq1_lenLoad[184] <= 32.0; sq1_lenLoad[185] <= 32.0; sq1_lenLoad[186] <= 32.0; sq1_lenLoad[187] <= 32.0; sq1_startVol[0] <= 12.0; sq1_startVol[1] <= 12.0; sq1_startVol[2] <= 12.0; sq1_startVol[3] <= 12.0; sq1_startVol[4] <= 12.0; sq1_startVol[5] <= 12.0; sq1_startVol[6] <= 12.0; sq1_startVol[7] <= 12.0; sq1_startVol[8] <= 12.0; sq1_startVol[9] <= 12.0; sq1_startVol[10] <= 12.0; sq1_startVol[11] <= 12.0; sq1_startVol[12] <= 12.0; sq1_startVol[13] <= 12.0; sq1_startVol[14] <= 12.0; sq1_startVol[15] <= 12.0; sq1_startVol[16] <= 12.0; sq1_startVol[17] <= 12.0; sq1_startVol[18] <= 12.0; sq1_startVol[19] <= 12.0; sq1_startVol[20] <= 12.0; sq1_startVol[21] <= 12.0; sq1_startVol[22] <= 12.0; sq1_startVol[23] <= 12.0; sq1_startVol[24] <= 12.0; sq1_startVol[25] <= 12.0; sq1_startVol[26] <= 12.0; sq1_startVol[27] <= 12.0; sq1_startVol[28] <= 12.0; sq1_startVol[29] <= 12.0; sq1_startVol[30] <= 12.0; sq1_startVol[31] <= 12.0; sq1_startVol[32] <= 12.0; sq1_startVol[33] <= 12.0; sq1_startVol[34] <= 12.0; sq1_startVol[35] <= 12.0; sq1_startVol[36] <= 12.0; sq1_startVol[37] <= 12.0; sq1_startVol[38] <= 12.0; sq1_startVol[39] <= 12.0; sq1_startVol[40] <= 12.0; sq1_startVol[41] <= 12.0; sq1_startVol[42] <= 12.0; sq1_startVol[43] <= 12.0; sq1_startVol[44] <= 12.0; sq1_startVol[45] <= 12.0; sq1_startVol[46] <= 12.0; sq1_startVol[47] <= 12.0; sq1_startVol[48] <= 12.0; sq1_startVol[49] <= 12.0; sq1_startVol[50] <= 12.0; sq1_startVol[51] <= 12.0; sq1_startVol[52] <= 12.0; sq1_startVol[53] <= 12.0; sq1_startVol[54] <= 12.0; sq1_startVol[55] <= 12.0; sq1_startVol[56] <= 12.0; sq1_startVol[57] <= 12.0; sq1_startVol[58] <= 12.0; sq1_startVol[59] <= 12.0; sq1_startVol[60] <= 12.0; sq1_startVol[61] <= 12.0; sq1_startVol[62] <= 12.0; sq1_startVol[63] <= 12.0; sq1_startVol[64] <= 12.0; sq1_startVol[65] <= 12.0; sq1_startVol[66] <= 12.0; sq1_startVol[67] <= 12.0; sq1_startVol[68] <= 12.0; sq1_startVol[69] <= 12.0; sq1_startVol[70] <= 12.0; sq1_startVol[71] <= 12.0; sq1_startVol[72] <= 12.0; sq1_startVol[73] <= 12.0; sq1_startVol[74] <= 12.0; sq1_startVol[75] <= 12.0; sq1_startVol[76] <= 12.0; sq1_startVol[77] <= 12.0; sq1_startVol[78] <= 12.0; sq1_startVol[79] <= 12.0; sq1_startVol[80] <= 12.0; sq1_startVol[81] <= 12.0; sq1_startVol[82] <= 12.0; sq1_startVol[83] <= 12.0; sq1_startVol[84] <= 12.0; sq1_startVol[85] <= 12.0; sq1_startVol[86] <= 12.0; sq1_startVol[87] <= 12.0; sq1_startVol[88] <= 12.0; sq1_startVol[89] <= 12.0; sq1_startVol[90] <= 12.0; sq1_startVol[91] <= 12.0; sq1_startVol[92] <= 12.0; sq1_startVol[93] <= 12.0; sq1_startVol[94] <= 12.0; sq1_startVol[95] <= 12.0; sq1_startVol[96] <= 12.0; sq1_startVol[97] <= 12.0; sq1_startVol[98] <= 12.0; sq1_startVol[99] <= 12.0; sq1_startVol[100] <= 12.0; sq1_startVol[101] <= 12.0; sq1_startVol[102] <= 12.0; sq1_startVol[103] <= 12.0; sq1_startVol[104] <= 12.0; sq1_startVol[105] <= 12.0; sq1_startVol[106] <= 12.0; sq1_startVol[107] <= 12.0; sq1_startVol[108] <= 12.0; sq1_startVol[109] <= 12.0; sq1_startVol[110] <= 12.0; sq1_startVol[111] <= 12.0; sq1_startVol[112] <= 12.0; sq1_startVol[113] <= 12.0; sq1_startVol[114] <= 12.0; sq1_startVol[115] <= 12.0; sq1_startVol[116] <= 12.0; sq1_startVol[117] <= 12.0; sq1_startVol[118] <= 12.0; sq1_startVol[119] <= 12.0; sq1_startVol[120] <= 12.0; sq1_startVol[121] <= 12.0; sq1_startVol[122] <= 12.0; sq1_startVol[123] <= 12.0; sq1_startVol[124] <= 12.0; sq1_startVol[125] <= 12.0; sq1_startVol[126] <= 12.0; sq1_startVol[127] <= 12.0; sq1_startVol[128] <= 12.0; sq1_startVol[129] <= 12.0; sq1_startVol[130] <= 12.0; sq1_startVol[131] <= 12.0; sq1_startVol[132] <= 12.0; sq1_startVol[133] <= 12.0; sq1_startVol[134] <= 12.0; sq1_startVol[135] <= 12.0; sq1_startVol[136] <= 12.0; sq1_startVol[137] <= 12.0; sq1_startVol[138] <= 12.0; sq1_startVol[139] <= 12.0; sq1_startVol[140] <= 12.0; sq1_startVol[141] <= 12.0; sq1_startVol[142] <= 12.0; sq1_startVol[143] <= 12.0; sq1_startVol[144] <= 12.0; sq1_startVol[145] <= 12.0; sq1_startVol[146] <= 12.0; sq1_startVol[147] <= 12.0; sq1_startVol[148] <= 12.0; sq1_startVol[149] <= 12.0; sq1_startVol[150] <= 12.0; sq1_startVol[151] <= 12.0; sq1_startVol[152] <= 12.0; sq1_startVol[153] <= 12.0; sq1_startVol[154] <= 12.0; sq1_startVol[155] <= 12.0; sq1_startVol[156] <= 12.0; sq1_startVol[157] <= 12.0; sq1_startVol[158] <= 12.0; sq1_startVol[159] <= 12.0; sq1_startVol[160] <= 12.0; sq1_startVol[161] <= 12.0; sq1_startVol[162] <= 12.0; sq1_startVol[163] <= 12.0; sq1_startVol[164] <= 12.0; sq1_startVol[165] <= 12.0; sq1_startVol[166] <= 12.0; sq1_startVol[167] <= 12.0; sq1_startVol[168] <= 12.0; sq1_startVol[169] <= 12.0; sq1_startVol[170] <= 12.0; sq1_startVol[171] <= 12.0; sq1_startVol[172] <= 12.0; sq1_startVol[173] <= 12.0; sq1_startVol[174] <= 12.0; sq1_startVol[175] <= 12.0; sq1_startVol[176] <= 12.0; sq1_startVol[177] <= 12.0; sq1_startVol[178] <= 12.0; sq1_startVol[179] <= 12.0; sq1_startVol[180] <= 12.0; sq1_startVol[181] <= 12.0; sq1_startVol[182] <= 12.0; sq1_startVol[183] <= 12.0; sq1_startVol[184] <= 12.0; sq1_startVol[185] <= 12.0; sq1_startVol[186] <= 12.0; sq1_startVol[187] <= 12.0; sq1_envAdd[0] <= 0.0; sq1_envAdd[1] <= 0.0; sq1_envAdd[2] <= 0.0; sq1_envAdd[3] <= 0.0; sq1_envAdd[4] <= 0.0; sq1_envAdd[5] <= 0.0; sq1_envAdd[6] <= 0.0; sq1_envAdd[7] <= 0.0; sq1_envAdd[8] <= 0.0; sq1_envAdd[9] <= 0.0; sq1_envAdd[10] <= 0.0; sq1_envAdd[11] <= 0.0; sq1_envAdd[12] <= 0.0; sq1_envAdd[13] <= 0.0; sq1_envAdd[14] <= 0.0; sq1_envAdd[15] <= 0.0; sq1_envAdd[16] <= 0.0; sq1_envAdd[17] <= 0.0; sq1_envAdd[18] <= 0.0; sq1_envAdd[19] <= 0.0; sq1_envAdd[20] <= 0.0; sq1_envAdd[21] <= 0.0; sq1_envAdd[22] <= 0.0; sq1_envAdd[23] <= 0.0; sq1_envAdd[24] <= 0.0; sq1_envAdd[25] <= 0.0; sq1_envAdd[26] <= 0.0; sq1_envAdd[27] <= 0.0; sq1_envAdd[28] <= 0.0; sq1_envAdd[29] <= 0.0; sq1_envAdd[30] <= 0.0; sq1_envAdd[31] <= 0.0; sq1_envAdd[32] <= 0.0; sq1_envAdd[33] <= 0.0; sq1_envAdd[34] <= 0.0; sq1_envAdd[35] <= 0.0; sq1_envAdd[36] <= 0.0; sq1_envAdd[37] <= 0.0; sq1_envAdd[38] <= 0.0; sq1_envAdd[39] <= 0.0; sq1_envAdd[40] <= 0.0; sq1_envAdd[41] <= 0.0; sq1_envAdd[42] <= 0.0; sq1_envAdd[43] <= 0.0; sq1_envAdd[44] <= 0.0; sq1_envAdd[45] <= 0.0; sq1_envAdd[46] <= 0.0; sq1_envAdd[47] <= 0.0; sq1_envAdd[48] <= 0.0; sq1_envAdd[49] <= 0.0; sq1_envAdd[50] <= 0.0; sq1_envAdd[51] <= 0.0; sq1_envAdd[52] <= 0.0; sq1_envAdd[53] <= 0.0; sq1_envAdd[54] <= 0.0; sq1_envAdd[55] <= 0.0; sq1_envAdd[56] <= 0.0; sq1_envAdd[57] <= 0.0; sq1_envAdd[58] <= 0.0; sq1_envAdd[59] <= 0.0; sq1_envAdd[60] <= 0.0; sq1_envAdd[61] <= 0.0; sq1_envAdd[62] <= 0.0; sq1_envAdd[63] <= 0.0; sq1_envAdd[64] <= 0.0; sq1_envAdd[65] <= 0.0; sq1_envAdd[66] <= 0.0; sq1_envAdd[67] <= 0.0; sq1_envAdd[68] <= 0.0; sq1_envAdd[69] <= 0.0; sq1_envAdd[70] <= 0.0; sq1_envAdd[71] <= 0.0; sq1_envAdd[72] <= 0.0; sq1_envAdd[73] <= 0.0; sq1_envAdd[74] <= 0.0; sq1_envAdd[75] <= 0.0; sq1_envAdd[76] <= 0.0; sq1_envAdd[77] <= 0.0; sq1_envAdd[78] <= 0.0; sq1_envAdd[79] <= 0.0; sq1_envAdd[80] <= 0.0; sq1_envAdd[81] <= 0.0; sq1_envAdd[82] <= 0.0; sq1_envAdd[83] <= 0.0; sq1_envAdd[84] <= 0.0; sq1_envAdd[85] <= 0.0; sq1_envAdd[86] <= 0.0; sq1_envAdd[87] <= 0.0; sq1_envAdd[88] <= 0.0; sq1_envAdd[89] <= 0.0; sq1_envAdd[90] <= 0.0; sq1_envAdd[91] <= 0.0; sq1_envAdd[92] <= 0.0; sq1_envAdd[93] <= 0.0; sq1_envAdd[94] <= 0.0; sq1_envAdd[95] <= 0.0; sq1_envAdd[96] <= 0.0; sq1_envAdd[97] <= 0.0; sq1_envAdd[98] <= 0.0; sq1_envAdd[99] <= 0.0; sq1_envAdd[100] <= 0.0; sq1_envAdd[101] <= 0.0; sq1_envAdd[102] <= 0.0; sq1_envAdd[103] <= 0.0; sq1_envAdd[104] <= 0.0; sq1_envAdd[105] <= 0.0; sq1_envAdd[106] <= 0.0; sq1_envAdd[107] <= 0.0; sq1_envAdd[108] <= 0.0; sq1_envAdd[109] <= 0.0; sq1_envAdd[110] <= 0.0; sq1_envAdd[111] <= 0.0; sq1_envAdd[112] <= 0.0; sq1_envAdd[113] <= 0.0; sq1_envAdd[114] <= 0.0; sq1_envAdd[115] <= 0.0; sq1_envAdd[116] <= 0.0; sq1_envAdd[117] <= 0.0; sq1_envAdd[118] <= 0.0; sq1_envAdd[119] <= 0.0; sq1_envAdd[120] <= 0.0; sq1_envAdd[121] <= 0.0; sq1_envAdd[122] <= 0.0; sq1_envAdd[123] <= 0.0; sq1_envAdd[124] <= 0.0; sq1_envAdd[125] <= 0.0; sq1_envAdd[126] <= 0.0; sq1_envAdd[127] <= 0.0; sq1_envAdd[128] <= 0.0; sq1_envAdd[129] <= 0.0; sq1_envAdd[130] <= 0.0; sq1_envAdd[131] <= 0.0; sq1_envAdd[132] <= 0.0; sq1_envAdd[133] <= 0.0; sq1_envAdd[134] <= 0.0; sq1_envAdd[135] <= 0.0; sq1_envAdd[136] <= 0.0; sq1_envAdd[137] <= 0.0; sq1_envAdd[138] <= 0.0; sq1_envAdd[139] <= 0.0; sq1_envAdd[140] <= 0.0; sq1_envAdd[141] <= 0.0; sq1_envAdd[142] <= 0.0; sq1_envAdd[143] <= 0.0; sq1_envAdd[144] <= 0.0; sq1_envAdd[145] <= 0.0; sq1_envAdd[146] <= 0.0; sq1_envAdd[147] <= 0.0; sq1_envAdd[148] <= 0.0; sq1_envAdd[149] <= 0.0; sq1_envAdd[150] <= 0.0; sq1_envAdd[151] <= 0.0; sq1_envAdd[152] <= 0.0; sq1_envAdd[153] <= 0.0; sq1_envAdd[154] <= 0.0; sq1_envAdd[155] <= 0.0; sq1_envAdd[156] <= 0.0; sq1_envAdd[157] <= 0.0; sq1_envAdd[158] <= 0.0; sq1_envAdd[159] <= 0.0; sq1_envAdd[160] <= 0.0; sq1_envAdd[161] <= 0.0; sq1_envAdd[162] <= 0.0; sq1_envAdd[163] <= 0.0; sq1_envAdd[164] <= 0.0; sq1_envAdd[165] <= 0.0; sq1_envAdd[166] <= 0.0; sq1_envAdd[167] <= 0.0; sq1_envAdd[168] <= 0.0; sq1_envAdd[169] <= 0.0; sq1_envAdd[170] <= 0.0; sq1_envAdd[171] <= 0.0; sq1_envAdd[172] <= 0.0; sq1_envAdd[173] <= 0.0; sq1_envAdd[174] <= 0.0; sq1_envAdd[175] <= 0.0; sq1_envAdd[176] <= 0.0; sq1_envAdd[177] <= 0.0; sq1_envAdd[178] <= 0.0; sq1_envAdd[179] <= 0.0; sq1_envAdd[180] <= 0.0; sq1_envAdd[181] <= 0.0; sq1_envAdd[182] <= 0.0; sq1_envAdd[183] <= 0.0; sq1_envAdd[184] <= 0.0; sq1_envAdd[185] <= 0.0; sq1_envAdd[186] <= 0.0; sq1_envAdd[187] <= 0.0; sq1_period[0] <= 4.0; sq1_period[1] <= 4.0; sq1_period[2] <= 4.0; sq1_period[3] <= 4.0; sq1_period[4] <= 4.0; sq1_period[5] <= 4.0; sq1_period[6] <= 4.0; sq1_period[7] <= 4.0; sq1_period[8] <= 4.0; sq1_period[9] <= 4.0; sq1_period[10] <= 4.0; sq1_period[11] <= 4.0; sq1_period[12] <= 4.0; sq1_period[13] <= 4.0; sq1_period[14] <= 4.0; sq1_period[15] <= 4.0; sq1_period[16] <= 4.0; sq1_period[17] <= 4.0; sq1_period[18] <= 4.0; sq1_period[19] <= 4.0; sq1_period[20] <= 4.0; sq1_period[21] <= 4.0; sq1_period[22] <= 4.0; sq1_period[23] <= 4.0; sq1_period[24] <= 4.0; sq1_period[25] <= 4.0; sq1_period[26] <= 4.0; sq1_period[27] <= 4.0; sq1_period[28] <= 4.0; sq1_period[29] <= 4.0; sq1_period[30] <= 4.0; sq1_period[31] <= 4.0; sq1_period[32] <= 4.0; sq1_period[33] <= 4.0; sq1_period[34] <= 4.0; sq1_period[35] <= 4.0; sq1_period[36] <= 4.0; sq1_period[37] <= 4.0; sq1_period[38] <= 4.0; sq1_period[39] <= 4.0; sq1_period[40] <= 4.0; sq1_period[41] <= 4.0; sq1_period[42] <= 4.0; sq1_period[43] <= 4.0; sq1_period[44] <= 4.0; sq1_period[45] <= 4.0; sq1_period[46] <= 4.0; sq1_period[47] <= 4.0; sq1_period[48] <= 4.0; sq1_period[49] <= 4.0; sq1_period[50] <= 4.0; sq1_period[51] <= 4.0; sq1_period[52] <= 4.0; sq1_period[53] <= 4.0; sq1_period[54] <= 4.0; sq1_period[55] <= 4.0; sq1_period[56] <= 4.0; sq1_period[57] <= 4.0; sq1_period[58] <= 4.0; sq1_period[59] <= 4.0; sq1_period[60] <= 4.0; sq1_period[61] <= 4.0; sq1_period[62] <= 4.0; sq1_period[63] <= 4.0; sq1_period[64] <= 4.0; sq1_period[65] <= 4.0; sq1_period[66] <= 4.0; sq1_period[67] <= 4.0; sq1_period[68] <= 4.0; sq1_period[69] <= 4.0; sq1_period[70] <= 4.0; sq1_period[71] <= 4.0; sq1_period[72] <= 4.0; sq1_period[73] <= 4.0; sq1_period[74] <= 4.0; sq1_period[75] <= 4.0; sq1_period[76] <= 4.0; sq1_period[77] <= 4.0; sq1_period[78] <= 4.0; sq1_period[79] <= 4.0; sq1_period[80] <= 4.0; sq1_period[81] <= 4.0; sq1_period[82] <= 4.0; sq1_period[83] <= 4.0; sq1_period[84] <= 4.0; sq1_period[85] <= 4.0; sq1_period[86] <= 4.0; sq1_period[87] <= 4.0; sq1_period[88] <= 4.0; sq1_period[89] <= 4.0; sq1_period[90] <= 4.0; sq1_period[91] <= 4.0; sq1_period[92] <= 4.0; sq1_period[93] <= 4.0; sq1_period[94] <= 4.0; sq1_period[95] <= 4.0; sq1_period[96] <= 4.0; sq1_period[97] <= 4.0; sq1_period[98] <= 4.0; sq1_period[99] <= 4.0; sq1_period[100] <= 4.0; sq1_period[101] <= 4.0; sq1_period[102] <= 4.0; sq1_period[103] <= 4.0; sq1_period[104] <= 4.0; sq1_period[105] <= 4.0; sq1_period[106] <= 4.0; sq1_period[107] <= 4.0; sq1_period[108] <= 4.0; sq1_period[109] <= 4.0; sq1_period[110] <= 4.0; sq1_period[111] <= 4.0; sq1_period[112] <= 4.0; sq1_period[113] <= 4.0; sq1_period[114] <= 4.0; sq1_period[115] <= 4.0; sq1_period[116] <= 4.0; sq1_period[117] <= 4.0; sq1_period[118] <= 4.0; sq1_period[119] <= 4.0; sq1_period[120] <= 4.0; sq1_period[121] <= 4.0; sq1_period[122] <= 4.0; sq1_period[123] <= 4.0; sq1_period[124] <= 4.0; sq1_period[125] <= 4.0; sq1_period[126] <= 4.0; sq1_period[127] <= 4.0; sq1_period[128] <= 4.0; sq1_period[129] <= 4.0; sq1_period[130] <= 4.0; sq1_period[131] <= 4.0; sq1_period[132] <= 4.0; sq1_period[133] <= 4.0; sq1_period[134] <= 4.0; sq1_period[135] <= 4.0; sq1_period[136] <= 4.0; sq1_period[137] <= 4.0; sq1_period[138] <= 4.0; sq1_period[139] <= 4.0; sq1_period[140] <= 4.0; sq1_period[141] <= 4.0; sq1_period[142] <= 4.0; sq1_period[143] <= 4.0; sq1_period[144] <= 4.0; sq1_period[145] <= 4.0; sq1_period[146] <= 4.0; sq1_period[147] <= 4.0; sq1_period[148] <= 4.0; sq1_period[149] <= 4.0; sq1_period[150] <= 4.0; sq1_period[151] <= 4.0; sq1_period[152] <= 4.0; sq1_period[153] <= 4.0; sq1_period[154] <= 4.0; sq1_period[155] <= 4.0; sq1_period[156] <= 4.0; sq1_period[157] <= 4.0; sq1_period[158] <= 4.0; sq1_period[159] <= 4.0; sq1_period[160] <= 4.0; sq1_period[161] <= 4.0; sq1_period[162] <= 4.0; sq1_period[163] <= 4.0; sq1_period[164] <= 4.0; sq1_period[165] <= 4.0; sq1_period[166] <= 4.0; sq1_period[167] <= 4.0; sq1_period[168] <= 4.0; sq1_period[169] <= 4.0; sq1_period[170] <= 4.0; sq1_period[171] <= 4.0; sq1_period[172] <= 4.0; sq1_period[173] <= 4.0; sq1_period[174] <= 4.0; sq1_period[175] <= 4.0; sq1_period[176] <= 4.0; sq1_period[177] <= 4.0; sq1_period[178] <= 4.0; sq1_period[179] <= 4.0; sq1_period[180] <= 4.0; sq1_period[181] <= 4.0; sq1_period[182] <= 4.0; sq1_period[183] <= 4.0; sq1_period[184] <= 4.0; sq1_period[185] <= 4.0; sq1_period[186] <= 4.0; sq1_period[187] <= 4.0; sq1_freq[0] <= 1546; sq1_freq[1] <= 1546; sq1_freq[2] <= 1546; sq1_freq[3] <= 1546; sq1_freq[4] <= 1546; sq1_freq[5] <= 1546; sq1_freq[6] <= 1546; sq1_freq[7] <= 1546; sq1_freq[8] <= 1602; sq1_freq[9] <= 1602; sq1_freq[10] <= 1602; sq1_freq[11] <= 1602; sq1_freq[12] <= 1602; sq1_freq[13] <= 1602; sq1_freq[14] <= 1602; sq1_freq[15] <= 1602; sq1_freq[16] <= 1546; sq1_freq[17] <= 1546; sq1_freq[18] <= 1546; sq1_freq[19] <= 1546; sq1_freq[20] <= 1546; sq1_freq[21] <= 1546; sq1_freq[22] <= 1546; sq1_freq[23] <= 1546; sq1_freq[24] <= 1673; sq1_freq[25] <= 1673; sq1_freq[26] <= 1673; sq1_freq[27] <= 1673; sq1_freq[28] <= 1673; sq1_freq[29] <= 1673; sq1_freq[30] <= 1673; sq1_freq[31] <= 1673; sq1_freq[32] <= 1650; sq1_freq[33] <= 1650; sq1_freq[34] <= 1650; sq1_freq[35] <= 1650; sq1_freq[36] <= 1650; sq1_freq[37] <= 1650; sq1_freq[38] <= 1650; sq1_freq[39] <= 1650; sq1_freq[40] <= 1650; sq1_freq[41] <= 1650; sq1_freq[42] <= 1650; sq1_freq[43] <= 1650; sq1_freq[44] <= 1650; sq1_freq[45] <= 1650; sq1_freq[46] <= 1650; sq1_freq[47] <= 1650; sq1_freq[48] <= 1546; sq1_freq[49] <= 1546; sq1_freq[50] <= 1546; sq1_freq[51] <= 1546; sq1_freq[52] <= 1546; sq1_freq[53] <= 1546; sq1_freq[54] <= 1546; sq1_freq[55] <= 1546; sq1_freq[56] <= 1602; sq1_freq[57] <= 1602; sq1_freq[58] <= 1602; sq1_freq[59] <= 1602; sq1_freq[60] <= 1602; sq1_freq[61] <= 1602; sq1_freq[62] <= 1602; sq1_freq[63] <= 1602; sq1_freq[64] <= 1546; sq1_freq[65] <= 1546; sq1_freq[66] <= 1546; sq1_freq[67] <= 1546; sq1_freq[68] <= 1546; sq1_freq[69] <= 1546; sq1_freq[70] <= 1546; sq1_freq[71] <= 1546; sq1_freq[72] <= 1714; sq1_freq[73] <= 1714; sq1_freq[74] <= 1714; sq1_freq[75] <= 1714; sq1_freq[76] <= 1714; sq1_freq[77] <= 1714; sq1_freq[78] <= 1714; sq1_freq[79] <= 1714; sq1_freq[80] <= 1673; sq1_freq[81] <= 1673; sq1_freq[82] <= 1673; sq1_freq[83] <= 1673; sq1_freq[84] <= 1673; sq1_freq[85] <= 1673; sq1_freq[86] <= 1673; sq1_freq[87] <= 1673; sq1_freq[88] <= 1673; sq1_freq[89] <= 1673; sq1_freq[90] <= 1673; sq1_freq[91] <= 1673; sq1_freq[92] <= 1673; sq1_freq[93] <= 1673; sq1_freq[94] <= 1673; sq1_freq[95] <= 1673; sq1_freq[96] <= 1546; sq1_freq[97] <= 1546; sq1_freq[98] <= 1546; sq1_freq[99] <= 1546; sq1_freq[100] <= 1546; sq1_freq[101] <= 1546; sq1_freq[102] <= 1546; sq1_freq[103] <= 1546; sq1_freq[104] <= 1798; sq1_freq[105] <= 1798; sq1_freq[106] <= 1798; sq1_freq[107] <= 1798; sq1_freq[108] <= 1798; sq1_freq[109] <= 1798; sq1_freq[110] <= 1798; sq1_freq[111] <= 1798; sq1_freq[112] <= 1750; sq1_freq[113] <= 1750; sq1_freq[114] <= 1750; sq1_freq[115] <= 1750; sq1_freq[116] <= 1750; sq1_freq[117] <= 1750; sq1_freq[118] <= 1750; sq1_freq[119] <= 1750; sq1_freq[120] <= 1673; sq1_freq[121] <= 1673; sq1_freq[122] <= 1673; sq1_freq[123] <= 1673; sq1_freq[124] <= 1673; sq1_freq[125] <= 1673; sq1_freq[126] <= 1673; sq1_freq[127] <= 1673; sq1_freq[128] <= 1650; sq1_freq[129] <= 1650; sq1_freq[130] <= 1650; sq1_freq[131] <= 1650; sq1_freq[132] <= 1650; sq1_freq[133] <= 1650; sq1_freq[134] <= 1650; sq1_freq[135] <= 1650; sq1_freq[136] <= 1602; sq1_freq[137] <= 1602; sq1_freq[138] <= 1602; sq1_freq[139] <= 1602; sq1_freq[140] <= 1602; sq1_freq[141] <= 1602; sq1_freq[142] <= 1602; sq1_freq[143] <= 1602; sq1_freq[144] <= 1602; sq1_freq[145] <= 1602; sq1_freq[146] <= 1602; sq1_freq[147] <= 1602; sq1_freq[148] <= 1602; sq1_freq[149] <= 1602; sq1_freq[150] <= 1602; sq1_freq[151] <= 1602; sq1_freq[152] <= 1767; sq1_freq[153] <= 1767; sq1_freq[154] <= 1767; sq1_freq[155] <= 1767; sq1_freq[156] <= 1767; sq1_freq[157] <= 1767; sq1_freq[158] <= 1767; sq1_freq[159] <= 1767; sq1_freq[160] <= 1750; sq1_freq[161] <= 1750; sq1_freq[162] <= 1750; sq1_freq[163] <= 1750; sq1_freq[164] <= 1750; sq1_freq[165] <= 1750; sq1_freq[166] <= 1750; sq1_freq[167] <= 1750; sq1_freq[168] <= 1673; sq1_freq[169] <= 1673; sq1_freq[170] <= 1673; sq1_freq[171] <= 1673; sq1_freq[172] <= 1673; sq1_freq[173] <= 1673; sq1_freq[174] <= 1673; sq1_freq[175] <= 1673; sq1_freq[176] <= 1714; sq1_freq[177] <= 1714; sq1_freq[178] <= 1714; sq1_freq[179] <= 1714; sq1_freq[180] <= 1714; sq1_freq[181] <= 1714; sq1_freq[182] <= 1714; sq1_freq[183] <= 1714; sq1_freq[184] <= 1673; sq1_freq[185] <= 1673; sq1_freq[186] <= 1673; sq1_freq[187] <= 1673; sq1_trigger[0] <= 1.0; sq1_trigger[1] <= 0; sq1_trigger[2] <= 0; sq1_trigger[3] <= 0; sq1_trigger[4] <= 0; sq1_trigger[5] <= 0; sq1_trigger[6] <= 1.0; sq1_trigger[7] <= 0; sq1_trigger[8] <= 1.0; sq1_trigger[9] <= 0; sq1_trigger[10] <= 0; sq1_trigger[11] <= 0; sq1_trigger[12] <= 0; sq1_trigger[13] <= 0; sq1_trigger[14] <= 0; sq1_trigger[15] <= 0; sq1_trigger[16] <= 1.0; sq1_trigger[17] <= 0; sq1_trigger[18] <= 0; sq1_trigger[19] <= 0; sq1_trigger[20] <= 0; sq1_trigger[21] <= 0; sq1_trigger[22] <= 0; sq1_trigger[23] <= 0; sq1_trigger[24] <= 1.0; sq1_trigger[25] <= 0; sq1_trigger[26] <= 0; sq1_trigger[27] <= 0; sq1_trigger[28] <= 0; sq1_trigger[29] <= 0; sq1_trigger[30] <= 0; sq1_trigger[31] <= 0; sq1_trigger[32] <= 1.0; sq1_trigger[33] <= 0; sq1_trigger[34] <= 0; sq1_trigger[35] <= 0; sq1_trigger[36] <= 0; sq1_trigger[37] <= 0; sq1_trigger[38] <= 0; sq1_trigger[39] <= 0; sq1_trigger[40] <= 0; sq1_trigger[41] <= 0; sq1_trigger[42] <= 0; sq1_trigger[43] <= 0; sq1_trigger[44] <= 0; sq1_trigger[45] <= 0; sq1_trigger[46] <= 0; sq1_trigger[47] <= 0; sq1_trigger[48] <= 1.0; sq1_trigger[49] <= 0; sq1_trigger[50] <= 0; sq1_trigger[51] <= 0; sq1_trigger[52] <= 0; sq1_trigger[53] <= 0; sq1_trigger[54] <= 1.0; sq1_trigger[55] <= 0; sq1_trigger[56] <= 1.0; sq1_trigger[57] <= 0; sq1_trigger[58] <= 0; sq1_trigger[59] <= 0; sq1_trigger[60] <= 0; sq1_trigger[61] <= 0; sq1_trigger[62] <= 0; sq1_trigger[63] <= 0; sq1_trigger[64] <= 1.0; sq1_trigger[65] <= 0; sq1_trigger[66] <= 0; sq1_trigger[67] <= 0; sq1_trigger[68] <= 0; sq1_trigger[69] <= 0; sq1_trigger[70] <= 0; sq1_trigger[71] <= 0; sq1_trigger[72] <= 1.0; sq1_trigger[73] <= 0; sq1_trigger[74] <= 0; sq1_trigger[75] <= 0; sq1_trigger[76] <= 0; sq1_trigger[77] <= 0; sq1_trigger[78] <= 0; sq1_trigger[79] <= 0; sq1_trigger[80] <= 1.0; sq1_trigger[81] <= 0; sq1_trigger[82] <= 0; sq1_trigger[83] <= 0; sq1_trigger[84] <= 0; sq1_trigger[85] <= 0; sq1_trigger[86] <= 0; sq1_trigger[87] <= 0; sq1_trigger[88] <= 0; sq1_trigger[89] <= 0; sq1_trigger[90] <= 0; sq1_trigger[91] <= 0; sq1_trigger[92] <= 0; sq1_trigger[93] <= 0; sq1_trigger[94] <= 0; sq1_trigger[95] <= 0; sq1_trigger[96] <= 1.0; sq1_trigger[97] <= 0; sq1_trigger[98] <= 0; sq1_trigger[99] <= 0; sq1_trigger[100] <= 0; sq1_trigger[101] <= 0; sq1_trigger[102] <= 1.0; sq1_trigger[103] <= 0; sq1_trigger[104] <= 1.0; sq1_trigger[105] <= 0; sq1_trigger[106] <= 0; sq1_trigger[107] <= 0; sq1_trigger[108] <= 0; sq1_trigger[109] <= 0; sq1_trigger[110] <= 0; sq1_trigger[111] <= 0; sq1_trigger[112] <= 1.0; sq1_trigger[113] <= 0; sq1_trigger[114] <= 0; sq1_trigger[115] <= 0; sq1_trigger[116] <= 0; sq1_trigger[117] <= 0; sq1_trigger[118] <= 0; sq1_trigger[119] <= 0; sq1_trigger[120] <= 1.0; sq1_trigger[121] <= 0; sq1_trigger[122] <= 0; sq1_trigger[123] <= 0; sq1_trigger[124] <= 0; sq1_trigger[125] <= 0; sq1_trigger[126] <= 0; sq1_trigger[127] <= 0; sq1_trigger[128] <= 1.0; sq1_trigger[129] <= 0; sq1_trigger[130] <= 0; sq1_trigger[131] <= 0; sq1_trigger[132] <= 0; sq1_trigger[133] <= 0; sq1_trigger[134] <= 0; sq1_trigger[135] <= 0; sq1_trigger[136] <= 1.0; sq1_trigger[137] <= 0; sq1_trigger[138] <= 0; sq1_trigger[139] <= 0; sq1_trigger[140] <= 0; sq1_trigger[141] <= 0; sq1_trigger[142] <= 0; sq1_trigger[143] <= 0; sq1_trigger[144] <= 0; sq1_trigger[145] <= 0; sq1_trigger[146] <= 0; sq1_trigger[147] <= 0; sq1_trigger[148] <= 0; sq1_trigger[149] <= 0; sq1_trigger[150] <= 0; sq1_trigger[151] <= 0; sq1_trigger[152] <= 1.0; sq1_trigger[153] <= 0; sq1_trigger[154] <= 0; sq1_trigger[155] <= 0; sq1_trigger[156] <= 0; sq1_trigger[157] <= 0; sq1_trigger[158] <= 1.0; sq1_trigger[159] <= 0; sq1_trigger[160] <= 1.0; sq1_trigger[161] <= 0; sq1_trigger[162] <= 0; sq1_trigger[163] <= 0; sq1_trigger[164] <= 0; sq1_trigger[165] <= 0; sq1_trigger[166] <= 0; sq1_trigger[167] <= 0; sq1_trigger[168] <= 1.0; sq1_trigger[169] <= 0; sq1_trigger[170] <= 0; sq1_trigger[171] <= 0; sq1_trigger[172] <= 0; sq1_trigger[173] <= 0; sq1_trigger[174] <= 0; sq1_trigger[175] <= 0; sq1_trigger[176] <= 1.0; sq1_trigger[177] <= 0; sq1_trigger[178] <= 0; sq1_trigger[179] <= 0; sq1_trigger[180] <= 0; sq1_trigger[181] <= 0; sq1_trigger[182] <= 0; sq1_trigger[183] <= 0; sq1_trigger[184] <= 1.0; sq1_trigger[185] <= 0; sq1_trigger[186] <= 0; sq1_trigger[187] <= 0; sq1_lenEnable[0] <= 1.0; sq1_lenEnable[1] <= 1.0; sq1_lenEnable[2] <= 1.0; sq1_lenEnable[3] <= 1.0; sq1_lenEnable[4] <= 1.0; sq1_lenEnable[5] <= 1.0; sq1_lenEnable[6] <= 1.0; sq1_lenEnable[7] <= 1.0; sq1_lenEnable[8] <= 1.0; sq1_lenEnable[9] <= 1.0; sq1_lenEnable[10] <= 1.0; sq1_lenEnable[11] <= 1.0; sq1_lenEnable[12] <= 1.0; sq1_lenEnable[13] <= 1.0; sq1_lenEnable[14] <= 1.0; sq1_lenEnable[15] <= 1.0; sq1_lenEnable[16] <= 1.0; sq1_lenEnable[17] <= 1.0; sq1_lenEnable[18] <= 1.0; sq1_lenEnable[19] <= 1.0; sq1_lenEnable[20] <= 1.0; sq1_lenEnable[21] <= 1.0; sq1_lenEnable[22] <= 1.0; sq1_lenEnable[23] <= 1.0; sq1_lenEnable[24] <= 1.0; sq1_lenEnable[25] <= 1.0; sq1_lenEnable[26] <= 1.0; sq1_lenEnable[27] <= 1.0; sq1_lenEnable[28] <= 1.0; sq1_lenEnable[29] <= 1.0; sq1_lenEnable[30] <= 1.0; sq1_lenEnable[31] <= 1.0; sq1_lenEnable[32] <= 1.0; sq1_lenEnable[33] <= 1.0; sq1_lenEnable[34] <= 1.0; sq1_lenEnable[35] <= 1.0; sq1_lenEnable[36] <= 1.0; sq1_lenEnable[37] <= 1.0; sq1_lenEnable[38] <= 1.0; sq1_lenEnable[39] <= 1.0; sq1_lenEnable[40] <= 1.0; sq1_lenEnable[41] <= 1.0; sq1_lenEnable[42] <= 1.0; sq1_lenEnable[43] <= 1.0; sq1_lenEnable[44] <= 1.0; sq1_lenEnable[45] <= 1.0; sq1_lenEnable[46] <= 1.0; sq1_lenEnable[47] <= 1.0; sq1_lenEnable[48] <= 1.0; sq1_lenEnable[49] <= 1.0; sq1_lenEnable[50] <= 1.0; sq1_lenEnable[51] <= 1.0; sq1_lenEnable[52] <= 1.0; sq1_lenEnable[53] <= 1.0; sq1_lenEnable[54] <= 1.0; sq1_lenEnable[55] <= 1.0; sq1_lenEnable[56] <= 1.0; sq1_lenEnable[57] <= 1.0; sq1_lenEnable[58] <= 1.0; sq1_lenEnable[59] <= 1.0; sq1_lenEnable[60] <= 1.0; sq1_lenEnable[61] <= 1.0; sq1_lenEnable[62] <= 1.0; sq1_lenEnable[63] <= 1.0; sq1_lenEnable[64] <= 1.0; sq1_lenEnable[65] <= 1.0; sq1_lenEnable[66] <= 1.0; sq1_lenEnable[67] <= 1.0; sq1_lenEnable[68] <= 1.0; sq1_lenEnable[69] <= 1.0; sq1_lenEnable[70] <= 1.0; sq1_lenEnable[71] <= 1.0; sq1_lenEnable[72] <= 1.0; sq1_lenEnable[73] <= 1.0; sq1_lenEnable[74] <= 1.0; sq1_lenEnable[75] <= 1.0; sq1_lenEnable[76] <= 1.0; sq1_lenEnable[77] <= 1.0; sq1_lenEnable[78] <= 1.0; sq1_lenEnable[79] <= 1.0; sq1_lenEnable[80] <= 1.0; sq1_lenEnable[81] <= 1.0; sq1_lenEnable[82] <= 1.0; sq1_lenEnable[83] <= 1.0; sq1_lenEnable[84] <= 1.0; sq1_lenEnable[85] <= 1.0; sq1_lenEnable[86] <= 1.0; sq1_lenEnable[87] <= 1.0; sq1_lenEnable[88] <= 1.0; sq1_lenEnable[89] <= 1.0; sq1_lenEnable[90] <= 1.0; sq1_lenEnable[91] <= 1.0; sq1_lenEnable[92] <= 1.0; sq1_lenEnable[93] <= 1.0; sq1_lenEnable[94] <= 1.0; sq1_lenEnable[95] <= 1.0; sq1_lenEnable[96] <= 1.0; sq1_lenEnable[97] <= 1.0; sq1_lenEnable[98] <= 1.0; sq1_lenEnable[99] <= 1.0; sq1_lenEnable[100] <= 1.0; sq1_lenEnable[101] <= 1.0; sq1_lenEnable[102] <= 1.0; sq1_lenEnable[103] <= 1.0; sq1_lenEnable[104] <= 1.0; sq1_lenEnable[105] <= 1.0; sq1_lenEnable[106] <= 1.0; sq1_lenEnable[107] <= 1.0; sq1_lenEnable[108] <= 1.0; sq1_lenEnable[109] <= 1.0; sq1_lenEnable[110] <= 1.0; sq1_lenEnable[111] <= 1.0; sq1_lenEnable[112] <= 1.0; sq1_lenEnable[113] <= 1.0; sq1_lenEnable[114] <= 1.0; sq1_lenEnable[115] <= 1.0; sq1_lenEnable[116] <= 1.0; sq1_lenEnable[117] <= 1.0; sq1_lenEnable[118] <= 1.0; sq1_lenEnable[119] <= 1.0; sq1_lenEnable[120] <= 1.0; sq1_lenEnable[121] <= 1.0; sq1_lenEnable[122] <= 1.0; sq1_lenEnable[123] <= 1.0; sq1_lenEnable[124] <= 1.0; sq1_lenEnable[125] <= 1.0; sq1_lenEnable[126] <= 1.0; sq1_lenEnable[127] <= 1.0; sq1_lenEnable[128] <= 1.0; sq1_lenEnable[129] <= 1.0; sq1_lenEnable[130] <= 1.0; sq1_lenEnable[131] <= 1.0; sq1_lenEnable[132] <= 1.0; sq1_lenEnable[133] <= 1.0; sq1_lenEnable[134] <= 1.0; sq1_lenEnable[135] <= 1.0; sq1_lenEnable[136] <= 1.0; sq1_lenEnable[137] <= 1.0; sq1_lenEnable[138] <= 1.0; sq1_lenEnable[139] <= 1.0; sq1_lenEnable[140] <= 1.0; sq1_lenEnable[141] <= 1.0; sq1_lenEnable[142] <= 1.0; sq1_lenEnable[143] <= 1.0; sq1_lenEnable[144] <= 1.0; sq1_lenEnable[145] <= 1.0; sq1_lenEnable[146] <= 1.0; sq1_lenEnable[147] <= 1.0; sq1_lenEnable[148] <= 1.0; sq1_lenEnable[149] <= 1.0; sq1_lenEnable[150] <= 1.0; sq1_lenEnable[151] <= 1.0; sq1_lenEnable[152] <= 1.0; sq1_lenEnable[153] <= 1.0; sq1_lenEnable[154] <= 1.0; sq1_lenEnable[155] <= 1.0; sq1_lenEnable[156] <= 1.0; sq1_lenEnable[157] <= 1.0; sq1_lenEnable[158] <= 1.0; sq1_lenEnable[159] <= 1.0; sq1_lenEnable[160] <= 1.0; sq1_lenEnable[161] <= 1.0; sq1_lenEnable[162] <= 1.0; sq1_lenEnable[163] <= 1.0; sq1_lenEnable[164] <= 1.0; sq1_lenEnable[165] <= 1.0; sq1_lenEnable[166] <= 1.0; sq1_lenEnable[167] <= 1.0; sq1_lenEnable[168] <= 1.0; sq1_lenEnable[169] <= 1.0; sq1_lenEnable[170] <= 1.0; sq1_lenEnable[171] <= 1.0; sq1_lenEnable[172] <= 1.0; sq1_lenEnable[173] <= 1.0; sq1_lenEnable[174] <= 1.0; sq1_lenEnable[175] <= 1.0; sq1_lenEnable[176] <= 1.0; sq1_lenEnable[177] <= 1.0; sq1_lenEnable[178] <= 1.0; sq1_lenEnable[179] <= 1.0; sq1_lenEnable[180] <= 1.0; sq1_lenEnable[181] <= 1.0; sq1_lenEnable[182] <= 1.0; sq1_lenEnable[183] <= 1.0; sq1_lenEnable[184] <= 1.0; sq1_lenEnable[185] <= 1.0; sq1_lenEnable[186] <= 1.0; sq1_lenEnable[187] <= 1.0;

	end

endmodule
